
module s38584 ( clk, rst, g35, g36, g6744, g6745, g6746, g6747, g6748, g6749, 
        g6750, g6751, g6752, g6753, g7243, g7245, g7257, g7260, g7540, g7916, 
        g7946, g8132, g8178, g8215, g8235, g8277, g8279, g8283, g8291, g8342, 
        g8344, g8353, g8358, g8398, g8403, g8416, g8475, g8719, g8783, g8784, 
        g8785, g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916, g8917, 
        g8918, g8919, g8920, g9019, g9048, g9251, g9497, g9553, g9555, g9615, 
        g9617, g9680, g9682, g9741, g9743, g9817, g10122, g10306, g10500, 
        g10527, g11349, g11388, g11418, g11447, g11678, g11770, g12184, g12238, 
        g12300, g12350, g12368, g12422, g12470, g12832, g12919, g12923, g13039, 
        g13049, g13068, g13085, g13099, g13259, g13272, g13865, g13881, g13895, 
        g13906, g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201, 
        g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673, g14694, 
        g14705, g14738, g14749, g14779, g14828, g16603, g16624, g16627, g16656, 
        g16659, g16686, g16693, g16718, g16722, g16744, g16748, g16775, g16874, 
        g16924, g16955, g17291, g17316, g17320, g17400, g17404, g17423, g17519, 
        g17577, g17580, g17604, g17607, g17639, g17646, g17649, g17674, g17678, 
        g17685, g17688, g17711, g17715, g17722, g17739, g17743, g17760, g17764, 
        g17778, g17787, g17813, g17819, g17845, g17871, g18092, g18094, g18095, 
        g18096, g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357, 
        g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176, g21245, 
        g21270, g21292, g21698, g21727, g23002, g23190, g23612, g23652, g23683, 
        g23759, g24151, g25114, g25167, g25219, g25259, g25582, g25583, g25584, 
        g25585, g25586, g25587, g25588, g25589, g25590, g26801, g26875, g26876, 
        g26877, g27831, g28030, g28041, g28042, g28753, g29210, g29211, g29212, 
        g29213, g29214, g29215, g29216, g29217, g29218, g29219, g29220, g29221, 
        g30327, g30329, g30330, g30331, g30332, g31521, g31656, g31665, g31793, 
        g31860, g31861, g31862, g31863, g32185, g32429, g32454, g32975, g33079, 
        g33435, g33533, g33636, g33659, g33874, g33894, g33935, g33945, g33946, 
        g33947, g33948, g33949, g33950, g33959, g34201, g34221, g34232, g34233, 
        g34234, g34235, g34236, g34237, g34238, g34239, g34240, g34383, g34425, 
        g34435, g34436, g34437, g34597, g34788, g34839, g34913, g34915, g34917, 
        g34919, g34921, g34923, g34925, g34927, g34956, g34972, test_se, 
        test_si );
  input clk, rst, g35, g36, g6744, g6745, g6746, g6747, g6748, g6749, g6750,
         g6751, g6752, g6753, test_se, test_si;
  output g7243, g7245, g7257, g7260, g7540, g7916, g7946, g8132, g8178, g8215,
         g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353, g8358, g8398,
         g8403, g8416, g8475, g8719, g8783, g8784, g8785, g8786, g8787, g8788,
         g8789, g8839, g8870, g8915, g8916, g8917, g8918, g8919, g8920, g9019,
         g9048, g9251, g9497, g9553, g9555, g9615, g9617, g9680, g9682, g9741,
         g9743, g9817, g10122, g10306, g10500, g10527, g11349, g11388, g11418,
         g11447, g11678, g11770, g12184, g12238, g12300, g12350, g12368,
         g12422, g12470, g12832, g12919, g12923, g13039, g13049, g13068,
         g13085, g13099, g13259, g13272, g13865, g13881, g13895, g13906,
         g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201,
         g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673,
         g14694, g14705, g14738, g14749, g14779, g14828, g16603, g16624,
         g16627, g16656, g16659, g16686, g16693, g16718, g16722, g16744,
         g16748, g16775, g16874, g16924, g16955, g17291, g17316, g17320,
         g17400, g17404, g17423, g17519, g17577, g17580, g17604, g17607,
         g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711,
         g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787,
         g17813, g17819, g17845, g17871, g18092, g18094, g18095, g18096,
         g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357,
         g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176,
         g21245, g21270, g21292, g21698, g21727, g23002, g23190, g23612,
         g23652, g23683, g23759, g24151, g25114, g25167, g25219, g25259,
         g25582, g25583, g25584, g25585, g25586, g25587, g25588, g25589,
         g25590, g26801, g26875, g26876, g26877, g27831, g28030, g28041,
         g28042, g28753, g29210, g29211, g29212, g29213, g29214, g29215,
         g29216, g29217, g29218, g29219, g29220, g29221, g30327, g30329,
         g30330, g30331, g30332, g31521, g31656, g31665, g31793, g31860,
         g31861, g31862, g31863, g32185, g32429, g32454, g32975, g33079,
         g33435, g33533, g33636, g33659, g33874, g33894, g33935, g33945,
         g33946, g33947, g33948, g33949, g33950, g33959, g34201, g34221,
         g34232, g34233, g34234, g34235, g34236, g34237, g34238, g34239,
         g34240, g34383, g34425, g34435, g34436, g34437, g34597, g34788,
         g34839, g34913, g34915, g34917, g34919, g34921, g34923, g34925,
         g34927, g34956, g34972;
  wire   g18092, g18094, g18095, g18096, g18097, g18098, g18099, g18100,
         g18101, g18881, g20049, g20557, g20652, g21176, g21245, g21270,
         g21292, g21698, g23002, g23652, g25114, g25167, g25219, g27831,
         g29211, g29212, g29215, g29219, g30329, g30331, g30332, g31862,
         g34435, g34788, g34956, g37, g4549, g4504, g2834, n716, n763, n4771,
         n4770, n4749, n7647, n721, n768, n671, n7805, n7809, n7596, n7813,
         n7618, n7817, n302, n7821, n7829, n7833, n7837, n3812, n3822, n3820,
         n3818, n3814, n3816, n3810, n7973, n7975, n7800, n603, n7825, n7826,
         n7824, n719, n699, n766, n7933, n7861, n7862, n7863, n7864, n7911,
         n7912, n7994, n7992, n7990, n489, n7986, n7984, n524, g26960, g4519,
         g4570, n7897, n7881, n7877, n5212, n5213, n5214, n5215, n5217, n5239,
         n5240, n5241, n5242, n5243, n5244, n5246, n5247, n5248, n5249, n5250,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5265,
         n5266, n5270, n5281, n5285, n5289, n5292, n5293, n5297, n5304, n5305,
         n5311, n5351, n5431, n5433, n5511, n5529, n5530, n5532, n5533, n5537,
         n5538, n5568, n5569, n5604, n5605, n5671, n5672, n5677, n5719, n5720,
         n5745, n5746, n5778, n5779, n5824, n5825, n5826, n5856, n5870, n5888,
         n5896, n5899, n5902, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6560, n6561, n6562, n6563, n6564, n6565,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n7045, n7046, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, g32975, g33959, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7801, n7802,
         n7803, n7804, n7806, n7807, n7808, n7810, n7811, n7812, n7814, n7815,
         n7816, n7818, n7819, n7820, n7822, n7823, n7827, n7828, n7830, n7831,
         n7832, n7834, n7835, n7836, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7878,
         n7879, n7880, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7974,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7985, n7987,
         n7988, n7989, n7991, n7993, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076;
  assign g34972 = 1'b1;
  assign g34927 = 1'b1;
  assign g34925 = 1'b1;
  assign g34923 = 1'b1;
  assign g34921 = 1'b1;
  assign g34919 = 1'b1;
  assign g34917 = 1'b1;
  assign g34915 = 1'b1;
  assign g34913 = 1'b1;
  assign g34437 = 1'b1;
  assign g34436 = 1'b1;
  assign g34425 = 1'b1;
  assign g34383 = 1'b1;
  assign g34240 = 1'b1;
  assign g34239 = 1'b1;
  assign g34238 = 1'b1;
  assign g34237 = 1'b1;
  assign g34236 = 1'b1;
  assign g34235 = 1'b1;
  assign g34234 = 1'b1;
  assign g34233 = 1'b1;
  assign g34232 = 1'b1;
  assign g34221 = 1'b1;
  assign g34201 = 1'b1;
  assign g33950 = 1'b1;
  assign g33949 = 1'b1;
  assign g33948 = 1'b1;
  assign g33947 = 1'b1;
  assign g33946 = 1'b1;
  assign g33945 = 1'b1;
  assign g33935 = 1'b1;
  assign g33874 = 1'b1;
  assign g33659 = 1'b1;
  assign g33636 = 1'b1;
  assign g32454 = 1'b1;
  assign g32429 = 1'b1;
  assign g31665 = 1'b1;
  assign g31656 = 1'b1;
  assign g25590 = 1'b1;
  assign g25589 = 1'b1;
  assign g25588 = 1'b1;
  assign g25587 = 1'b1;
  assign g25586 = 1'b1;
  assign g25585 = 1'b1;
  assign g25584 = 1'b1;
  assign g25583 = 1'b1;
  assign g25582 = 1'b1;
  assign g24151 = 1'b1;
  assign g23190 = 1'b1;
  assign g34597 = 1'b0;
  assign g12368 = 1'b0;
  assign g9048 = 1'b0;
  assign g8403 = 1'b0;
  assign g8353 = 1'b0;
  assign g8283 = 1'b0;
  assign g8235 = 1'b0;
  assign g8178 = 1'b0;
  assign g8132 = 1'b0;
  assign g18092 = g6753;
  assign g18094 = g6748;
  assign g18095 = g6749;
  assign g18096 = g6750;
  assign g18097 = g6747;
  assign g18098 = g6744;
  assign g18099 = g6745;
  assign g18100 = g6751;
  assign g18101 = g6746;
  assign g29218 = g18881;
  assign g29210 = g20049;
  assign g29213 = g20557;
  assign g29214 = g20652;
  assign g29216 = g21176;
  assign g29220 = g21245;
  assign g29217 = g21270;
  assign g29221 = g21292;
  assign g21698 = g36;
  assign g30327 = g23002;
  assign g30330 = g23652;
  assign g31860 = g25114;
  assign g31863 = g25167;
  assign g31861 = g25219;
  assign g33533 = g27831;
  assign g20763 = g29211;
  assign g20899 = g29212;
  assign g20901 = g29215;
  assign g20654 = g29219;
  assign g23612 = g30329;
  assign g23759 = g30331;
  assign g23683 = g30332;
  assign g25259 = g31862;
  assign g31521 = g34435;
  assign g33894 = g34788;
  assign g34839 = g34956;
  assign g26801 = g32975;
  assign g28753 = g33959;

  DFFSRX1 g859_reg ( .D(n7063), .CK(clk), .RN(n7987), .SN(1'b1), .Q(g14189), 
        .QN(n5899) );
  DFFSRX1 g869_reg ( .D(n7070), .CK(clk), .RN(n7985), .SN(1'b1), .Q(g14201) );
  DFFSRX1 g875_reg ( .D(n7068), .CK(clk), .RN(n8085), .SN(1'b1), .Q(g14217) );
  DFFSRX1 g878_reg ( .D(g14217), .CK(clk), .RN(n8085), .SN(1'b1), .Q(g14096)
         );
  DFFSRX1 g881_reg ( .D(g14096), .CK(clk), .RN(n8085), .SN(1'b1), .Q(g14125)
         );
  DFFSRX1 g884_reg ( .D(g14125), .CK(clk), .RN(n8085), .SN(1'b1), .Q(g14147)
         );
  DFFSRX1 g887_reg ( .D(g14147), .CK(clk), .RN(n8085), .SN(1'b1), .Q(g14167), 
        .QN(n5896) );
  DFFSRX1 g872_reg ( .D(n7069), .CK(clk), .RN(n8085), .SN(1'b1), .Q(n12772) );
  DFFSRX1 g2084_reg ( .D(n7122), .CK(clk), .RN(n8000), .SN(1'b1), .Q(n12799)
         );
  DFFSRX1 g2241_reg ( .D(n7123), .CK(clk), .RN(n7989), .SN(1'b1), .Q(n12776)
         );
  DFFSRX1 g2852_reg ( .D(n7139), .CK(clk), .RN(n8080), .SN(1'b1), .Q(n12682), 
        .QN(n7770) );
  DFFSRX1 g2856_reg ( .D(n7163), .CK(clk), .RN(n7988), .SN(1'b1), .Q(n12681), 
        .QN(n7740) );
  DFFSRX1 g2860_reg ( .D(n7140), .CK(clk), .RN(n8080), .SN(1'b1), .Q(n12680), 
        .QN(n7785) );
  DFFSRX1 g2932_reg ( .D(n7202), .CK(clk), .RN(n8058), .SN(1'b1), .Q(n12650), 
        .QN(n7834) );
  DFFSRX1 g2984_reg ( .D(n7049), .CK(clk), .RN(n8079), .SN(1'b1), .Q(n12657), 
        .QN(n7743) );
  DFFSRX1 g2994_reg ( .D(n7142), .CK(clk), .RN(n7985), .SN(1'b1), .Q(n12640), 
        .QN(n7768) );
  DFFSRX1 g2999_reg ( .D(n7173), .CK(clk), .RN(n7985), .SN(1'b1), .Q(n12639)
         );
  DFFSRX1 g3050_reg ( .D(n7155), .CK(clk), .RN(n8081), .SN(1'b1), .Q(n12638)
         );
  DFFSRX1 g3100_reg ( .D(n7094), .CK(clk), .RN(n8081), .SN(1'b1), .Q(n12637), 
        .QN(n7776) );
  DFFSRX1 g3147_reg ( .D(n7099), .CK(clk), .RN(n8069), .SN(1'b1), .Q(n12599), 
        .QN(n7745) );
  DFFSRX1 g3111_reg ( .D(n7109), .CK(clk), .RN(n8068), .SN(1'b1), .Q(n12634), 
        .QN(n7675) );
  DFFSRX1 g4944_reg ( .D(n7062), .CK(clk), .RN(n8067), .SN(1'b1), .Q(n12550), 
        .QN(n7698) );
  DFFSRX1 g4950_reg ( .D(n7171), .CK(clk), .RN(n8032), .SN(1'b1), .Q(n12301), 
        .QN(n7778) );
  DFFSRX1 g4955_reg ( .D(n7133), .CK(clk), .RN(n8032), .SN(1'b1), .Q(n12523), 
        .QN(n7704) );
  DFFSRX1 g4961_reg ( .D(n7107), .CK(clk), .RN(n8037), .SN(1'b1), .Q(n12300), 
        .QN(n7789) );
  DFFSRX1 g4572_reg ( .D(n7046), .CK(clk), .RN(n8078), .SN(1'b1), .Q(n12393)
         );
  DFFSRX1 g4575_reg ( .D(n7177), .CK(clk), .RN(n7988), .SN(1'b1), .Q(n12406)
         );
  DFFSRX1 g4578_reg ( .D(n7178), .CK(clk), .RN(n7988), .SN(1'b1), .Q(n12386), 
        .QN(n7836) );
  DFFSRX1 g5503_reg ( .D(n7103), .CK(clk), .RN(n8043), .SN(1'b1), .Q(n12235)
         );
  DFFSRX1 g5467_reg ( .D(n7113), .CK(clk), .RN(n8042), .SN(1'b1), .Q(n12238), 
        .QN(n7710) );
  DFFSRX1 g5673_reg ( .D(n7078), .CK(clk), .RN(n8039), .SN(1'b1), .Q(g17813), 
        .QN(n5259) );
  DFFSRX1 g5677_reg ( .D(g17813), .CK(clk), .RN(n8039), .SN(1'b1), .Q(g14635), 
        .QN(n5258) );
  DFFSRX1 g4821_reg ( .D(n7128), .CK(clk), .RN(n8039), .SN(1'b1), .Q(n12394), 
        .QN(n7783) );
  DFFSRX1 g4831_reg ( .D(n7129), .CK(clk), .RN(n8069), .SN(1'b1), .Q(n12396)
         );
  DFFSRX1 g3317_reg ( .D(n7093), .CK(clk), .RN(n8048), .SN(1'b1), .Q(g16874)
         );
  DFFSRX1 g3321_reg ( .D(g16874), .CK(clk), .RN(n8048), .SN(1'b1), .Q(g13865)
         );
  DFFSRX1 g3401_reg ( .D(n7156), .CK(clk), .RN(n8065), .SN(1'b1), .Q(n12584)
         );
  DFFSRX1 g3451_reg ( .D(n7092), .CK(clk), .RN(n8065), .SN(1'b1), .Q(n12583), 
        .QN(n7775) );
  DFFSRX1 g3498_reg ( .D(n7100), .CK(clk), .RN(n8066), .SN(1'b1), .Q(n12545)
         );
  DFFSRX1 g3462_reg ( .D(n7110), .CK(clk), .RN(n8064), .SN(1'b1), .Q(n12548)
         );
  DFFSRX1 g3684_reg ( .D(n7127), .CK(clk), .RN(n8065), .SN(1'b1), .Q(n12531)
         );
  DFFSRX1 g3752_reg ( .D(n7157), .CK(clk), .RN(n8064), .SN(1'b1), .Q(n12528)
         );
  DFFSRX1 g3802_reg ( .D(n7090), .CK(clk), .RN(n8063), .SN(1'b1), .Q(n12527), 
        .QN(n7748) );
  DFFSRX1 g3849_reg ( .D(n7101), .CK(clk), .RN(n8063), .SN(1'b1), .Q(n12497)
         );
  DFFSRX1 g3813_reg ( .D(n7111), .CK(clk), .RN(n8063), .SN(1'b1), .Q(n12500), 
        .QN(n7711) );
  DFFSRX1 g4157_reg ( .D(n7143), .CK(clk), .RN(n8060), .SN(1'b1), .Q(n12471)
         );
  DFFSRX1 g4191_reg ( .D(n7182), .CK(clk), .RN(n8060), .SN(1'b1), .Q(g11447), 
        .QN(n5243) );
  DFFSRX1 g4194_reg ( .D(n7087), .CK(clk), .RN(n8059), .SN(1'b1), .Q(g8784), 
        .QN(n5241) );
  DFFSRX1 g4200_reg ( .D(g8785), .CK(clk), .RN(n8059), .SN(1'b1), .Q(g8786), 
        .QN(n5240) );
  DFFSRX1 g4219_reg ( .D(g8916), .CK(clk), .RN(n8059), .SN(1'b1), .Q(g8917), 
        .QN(n5217) );
  DFFSRX1 g4226_reg ( .D(g8870), .CK(clk), .RN(n8059), .SN(1'b1), .Q(g8918), 
        .QN(n5215) );
  DFFSRX1 g4229_reg ( .D(g8918), .CK(clk), .RN(n8059), .SN(1'b1), .Q(g8919), 
        .QN(n5214) );
  DFFSRX1 g4232_reg ( .D(g8919), .CK(clk), .RN(n8058), .SN(1'b1), .Q(g8920), 
        .QN(n5213) );
  DFFSRX1 g4245_reg ( .D(n7154), .CK(clk), .RN(n8058), .SN(1'b1), .Q(n12465), 
        .QN(n7777) );
  DFFSRX1 g4249_reg ( .D(n7144), .CK(clk), .RN(n8058), .SN(1'b1), .Q(n12464), 
        .QN(n7794) );
  DFFSRX1 g4188_reg ( .D(n7088), .CK(clk), .RN(n8037), .SN(1'b1), .Q(g8783), 
        .QN(n5242) );
  DFFSRX1 g4258_reg ( .D(n7057), .CK(clk), .RN(n8058), .SN(1'b1), .Q(n12460), 
        .QN(n7625) );
  DFFSRX1 g4277_reg ( .D(n7183), .CK(clk), .RN(n8057), .SN(1'b1), .Q(g8839), 
        .QN(n5244) );
  DFFSRX1 g4284_reg ( .D(n7058), .CK(clk), .RN(n8057), .SN(1'b1), .Q(n12593)
         );
  DFFSRX1 g4287_reg ( .D(n7051), .CK(clk), .RN(n8057), .SN(1'b1), .Q(g9019), 
        .QN(n5856) );
  DFFSRX1 g4297_reg ( .D(g10122), .CK(clk), .RN(n8037), .SN(1'b1), .Q(n12458)
         );
  DFFSRX1 g4304_reg ( .D(n7059), .CK(clk), .RN(n8058), .SN(1'b1), .Q(g9251), 
        .QN(n5212) );
  DFFSRX1 g4308_reg ( .D(g9251), .CK(clk), .RN(n8058), .SN(1'b1), .Q(n12653), 
        .QN(n7623) );
  DFFSRX1 g4366_reg ( .D(n7060), .CK(clk), .RN(n7988), .SN(1'b1), .Q(n12538), 
        .QN(n7762) );
  DFFSRX1 g4019_reg ( .D(n7089), .CK(clk), .RN(n8031), .SN(1'b1), .Q(g16955), 
        .QN(n5248) );
  DFFSRX1 g4023_reg ( .D(g16955), .CK(clk), .RN(n8031), .SN(1'b1), .Q(g13906), 
        .QN(n5247) );
  DFFSRX1 g3668_reg ( .D(n7091), .CK(clk), .RN(n8064), .SN(1'b1), .Q(g16924), 
        .QN(n5250) );
  DFFSRX1 g3672_reg ( .D(g16924), .CK(clk), .RN(n8064), .SN(1'b1), .Q(g13881), 
        .QN(n5249) );
  DFFSRX1 g6541_reg ( .D(n7098), .CK(clk), .RN(n8036), .SN(1'b1), .Q(n12180)
         );
  DFFSRX1 g5011_reg ( .D(n7130), .CK(clk), .RN(n8034), .SN(1'b1), .Q(n12387)
         );
  DFFSRX1 g5109_reg ( .D(n7082), .CK(clk), .RN(n8029), .SN(1'b1), .Q(n12266), 
        .QN(n7797) );
  DFFSRX1 g5112_reg ( .D(n7081), .CK(clk), .RN(n8029), .SN(1'b1), .Q(n12272), 
        .QN(n7774) );
  DFFSRX1 g5022_reg ( .D(n7158), .CK(clk), .RN(n8029), .SN(1'b1), .Q(n12278)
         );
  DFFSRX1 g5156_reg ( .D(n7102), .CK(clk), .RN(n8074), .SN(1'b1), .Q(n12254)
         );
  DFFSRX1 g5120_reg ( .D(n7112), .CK(clk), .RN(n8028), .SN(1'b1), .Q(n12258), 
        .QN(n7713) );
  DFFSRX1 g5327_reg ( .D(n7080), .CK(clk), .RN(n8072), .SN(1'b1), .Q(g17787), 
        .QN(n5261) );
  DFFSRX1 g5331_reg ( .D(g17787), .CK(clk), .RN(n8072), .SN(1'b1), .Q(g14597), 
        .QN(n5260) );
  DFFSRX1 g5406_reg ( .D(n7159), .CK(clk), .RN(n8040), .SN(1'b1), .Q(n12244)
         );
  DFFSRX1 g5456_reg ( .D(n7079), .CK(clk), .RN(n8040), .SN(1'b1), .Q(n12243), 
        .QN(n7747) );
  DFFSRX1 g4754_reg ( .D(n7061), .CK(clk), .RN(n8071), .SN(1'b1), .Q(n12402), 
        .QN(n7699) );
  DFFSRX1 g4760_reg ( .D(n7169), .CK(clk), .RN(n8044), .SN(1'b1), .Q(n12379), 
        .QN(n7669) );
  DFFSRX1 g4765_reg ( .D(n7131), .CK(clk), .RN(n8044), .SN(1'b1), .Q(n12400), 
        .QN(n7701) );
  DFFSRX1 g4771_reg ( .D(n7165), .CK(clk), .RN(n8045), .SN(1'b1), .Q(n12375), 
        .QN(n7801) );
  DFFSRX1 g5817_reg ( .D(n7164), .CK(clk), .RN(n8071), .SN(1'b1), .Q(n12679), 
        .QN(n7331) );
  DFFSRX1 g5849_reg ( .D(n7104), .CK(clk), .RN(n8070), .SN(1'b1), .Q(n12209)
         );
  DFFSRX1 g5813_reg ( .D(n7114), .CK(clk), .RN(n8030), .SN(1'b1), .Q(n12213), 
        .QN(n7702) );
  DFFSRX1 g6019_reg ( .D(n7076), .CK(clk), .RN(n8052), .SN(1'b1), .Q(g17819), 
        .QN(n5257) );
  DFFSRX1 g6023_reg ( .D(g17819), .CK(clk), .RN(n8052), .SN(1'b1), .Q(g14673), 
        .QN(n5256) );
  DFFSRX1 g5802_reg ( .D(n7077), .CK(clk), .RN(n8040), .SN(1'b1), .Q(n12215), 
        .QN(n7773) );
  DFFSRX1 g5752_reg ( .D(n7160), .CK(clk), .RN(n8040), .SN(1'b1), .Q(n12216)
         );
  DFFSRX1 g6163_reg ( .D(n7153), .CK(clk), .RN(n8038), .SN(1'b1), .Q(n12677), 
        .QN(n7621) );
  DFFSRX1 g6195_reg ( .D(n7105), .CK(clk), .RN(n8048), .SN(1'b1), .Q(n12195)
         );
  DFFSRX1 g6159_reg ( .D(n7115), .CK(clk), .RN(n8038), .SN(1'b1), .Q(n12199), 
        .QN(n7668) );
  DFFSRX1 g6365_reg ( .D(n7074), .CK(clk), .RN(n8044), .SN(1'b1), .Q(g17845), 
        .QN(n5255) );
  DFFSRX1 g6369_reg ( .D(g17845), .CK(clk), .RN(n8044), .SN(1'b1), .Q(g14705), 
        .QN(n5254) );
  DFFSRX1 g6148_reg ( .D(n7075), .CK(clk), .RN(n8038), .SN(1'b1), .Q(n12201), 
        .QN(n7772) );
  DFFSRX1 g6098_reg ( .D(n7161), .CK(clk), .RN(n8038), .SN(1'b1), .Q(n12202)
         );
  DFFSRX1 g94_reg ( .D(n7191), .CK(clk), .RN(n8025), .SN(1'b1), .Q(g20652), 
        .QN(n5870) );
  DFFSRX1 g102_reg ( .D(n7198), .CK(clk), .RN(n8026), .SN(1'b1), .Q(g29215) );
  DFFSRX1 g1075_reg ( .D(n7194), .CK(clk), .RN(n8021), .SN(1'b1), .Q(g17291), 
        .QN(n5246) );
  DFFSRX1 g1087_reg ( .D(g17400), .CK(clk), .RN(n8021), .SN(1'b1), .Q(n13048)
         );
  DFFSRX1 g1111_reg ( .D(n7167), .CK(clk), .RN(n8022), .SN(1'b1), .Q(n13039)
         );
  DFFSRX1 g1141_reg ( .D(n7117), .CK(clk), .RN(n8022), .SN(1'b1), .Q(n13034), 
        .QN(n7611) );
  DFFSRX1 g496_reg ( .D(n7197), .CK(clk), .RN(n8025), .SN(1'b1), .Q(n12896) );
  DFFSRX1 g1418_reg ( .D(n7195), .CK(clk), .RN(n8018), .SN(1'b1), .Q(g17320), 
        .QN(n5266) );
  DFFSRX1 g1484_reg ( .D(n7118), .CK(clk), .RN(n8014), .SN(1'b1), .Q(n12970), 
        .QN(n7717) );
  DFFSRX1 g1454_reg ( .D(n7168), .CK(clk), .RN(n8017), .SN(1'b1), .Q(n12910)
         );
  DFFSRX1 g79_reg ( .D(n7199), .CK(clk), .RN(n8025), .SN(1'b1), .Q(g29212), 
        .QN(n5533) );
  DFFSRX1 g686_reg ( .D(n7116), .CK(clk), .RN(n8083), .SN(1'b1), .Q(n12328) );
  DFFSRX1 g728_reg ( .D(n7170), .CK(clk), .RN(n8025), .SN(1'b1), .Q(n12169) );
  DFFSRX1 g736_reg ( .D(n7071), .CK(clk), .RN(n8085), .SN(1'b1), .Q(n12241) );
  DFFSRX1 g799_reg ( .D(n7067), .CK(clk), .RN(n8085), .SN(1'b1), .Q(g12184) );
  DFFSRX1 g355_reg ( .D(n7050), .CK(clk), .RN(n8027), .SN(1'b1), .Q(n12532), 
        .QN(n7705) );
  DFFSRX1 g365_reg ( .D(n7201), .CK(clk), .RN(n8027), .SN(1'b1), .Q(g8719), 
        .QN(n5902) );
  DFFSRX1 g429_reg ( .D(n7097), .CK(clk), .RN(n8023), .SN(1'b1), .Q(n12487) );
  DFFSRX1 g203_reg ( .D(n7200), .CK(clk), .RN(n8012), .SN(1'b1), .Q(n12906), 
        .QN(n7841) );
  DFFSRX1 g215_reg ( .D(n7048), .CK(clk), .RN(n8011), .SN(1'b1), .Q(g8291), 
        .QN(n7828) );
  DFFSRX1 g222_reg ( .D(n7196), .CK(clk), .RN(n8012), .SN(1'b1), .Q(n12827) );
  DFFSRX1 g433_reg ( .D(n7108), .CK(clk), .RN(n8023), .SN(1'b1), .Q(n12457), 
        .QN(n7812) );
  DFFSRX1 g504_reg ( .D(n7106), .CK(clk), .RN(n8025), .SN(1'b1), .Q(n12267) );
  DFFSRX1 g538_reg ( .D(n7174), .CK(clk), .RN(n8012), .SN(1'b1), .Q(n12245), 
        .QN(n7810) );
  DFFSRX1 g117_reg ( .D(n7180), .CK(clk), .RN(n7997), .SN(1'b1), .Q(g21270), 
        .QN(n5265) );
  DFFSRX1 g121_reg ( .D(n7181), .CK(clk), .RN(n7997), .SN(1'b1), .Q(g29219) );
  DFFSRX1 g2204_reg ( .D(n7135), .CK(clk), .RN(n7989), .SN(1'b1), .Q(n12779), 
        .QN(n7693) );
  DFFSRX1 g2223_reg ( .D(n7150), .CK(clk), .RN(n7991), .SN(1'b1), .Q(n12778), 
        .QN(n7234) );
  DFFSRX1 g2375_reg ( .D(n7124), .CK(clk), .RN(n8010), .SN(1'b1), .Q(n12749)
         );
  DFFSRX1 g2338_reg ( .D(n7151), .CK(clk), .RN(n7991), .SN(1'b1), .Q(n12751), 
        .QN(n7347) );
  DFFSRX1 g2357_reg ( .D(n7152), .CK(clk), .RN(n7993), .SN(1'b1), .Q(n12750), 
        .QN(n7210) );
  DFFSRX1 g2509_reg ( .D(n7125), .CK(clk), .RN(n8010), .SN(1'b1), .Q(n12728)
         );
  DFFSRX1 g2472_reg ( .D(n7136), .CK(clk), .RN(n7998), .SN(1'b1), .Q(n12730), 
        .QN(n7694) );
  DFFSRX1 g2643_reg ( .D(n7126), .CK(clk), .RN(n7996), .SN(1'b1), .Q(n12707)
         );
  DFFSRX1 g2606_reg ( .D(n7137), .CK(clk), .RN(n7996), .SN(1'b1), .Q(n12709), 
        .QN(n7348) );
  DFFSRX1 g2763_reg ( .D(n7193), .CK(clk), .RN(n8007), .SN(1'b1), .QN(n5351)
         );
  DFFSRX1 g1682_reg ( .D(n7119), .CK(clk), .RN(n8005), .SN(1'b1), .Q(n12875)
         );
  DFFSRX1 g1644_reg ( .D(n7145), .CK(clk), .RN(n8004), .SN(1'b1), .Q(n12877), 
        .QN(n7691) );
  DFFSRX1 g1664_reg ( .D(n7146), .CK(clk), .RN(n8003), .SN(1'b1), .Q(n12876), 
        .QN(n7232) );
  DFFSRX1 g1816_reg ( .D(n7120), .CK(clk), .RN(n8002), .SN(1'b1), .Q(n12853)
         );
  DFFSRX1 g1779_reg ( .D(n7147), .CK(clk), .RN(n8001), .SN(1'b1), .Q(n12855), 
        .QN(n7345) );
  DFFSRX1 g1798_reg ( .D(n7148), .CK(clk), .RN(n8001), .SN(1'b1), .Q(n12854), 
        .QN(n7208) );
  DFFSRX1 g1950_reg ( .D(n7121), .CK(clk), .RN(n8006), .SN(1'b1), .Q(n12826), 
        .QN(n7703) );
  DFFSRX1 g1913_reg ( .D(n7134), .CK(clk), .RN(n7998), .SN(1'b1), .Q(n12831), 
        .QN(n7692) );
  DFFSRX1 g1932_reg ( .D(n7149), .CK(clk), .RN(n8007), .SN(1'b1), .Q(n12830), 
        .QN(n7233) );
  DFFSRX1 g2878_reg ( .D(n7179), .CK(clk), .RN(n7985), .SN(1'b1), .Q(n12664), 
        .QN(n7842) );
  DFFSRX1 g2890_reg ( .D(n7184), .CK(clk), .RN(n8080), .SN(1'b1), .Q(n12684), 
        .QN(n7832) );
  DFFSRX1 g2894_reg ( .D(n7141), .CK(clk), .RN(n8080), .SN(1'b1), .Q(n12661), 
        .QN(n7786) );
  DFFSRX1 g59_reg ( .D(n7045), .CK(clk), .RN(n7988), .SN(1'b1), .Q(g20049), 
        .QN(n5239) );
  DFFSRX1 g66_reg ( .D(n7192), .CK(clk), .RN(n8027), .SN(1'b1), .Q(g18881) );
  DFFSRX1 g4537_reg ( .D(n7187), .CK(clk), .RN(n8079), .SN(1'b1), .Q(g10306), 
        .QN(n5311) );
  DFFSRX1 g4430_reg ( .D(n7172), .CK(clk), .RN(n7987), .SN(1'b1), .Q(n12433), 
        .QN(n7815) );
  DFFSRX1 g4455_reg ( .D(n7086), .CK(clk), .RN(n8076), .SN(1'b1), .Q(n12812)
         );
  DFFSRX1 g4456_reg ( .D(n7066), .CK(clk), .RN(n8076), .SN(1'b1), .Q(n12426), 
        .QN(n7843) );
  DFFSRX1 g4474_reg ( .D(n7085), .CK(clk), .RN(n8076), .SN(1'b1), .Q(g26960)
         );
  DFFSRX1 g4477_reg ( .D(g26960), .CK(clk), .RN(n8076), .SN(1'b1), .QN(n5297)
         );
  DFFSRX1 g4483_reg ( .D(n7084), .CK(clk), .RN(n7987), .SN(1'b1), .Q(n12419)
         );
  DFFSRX1 g4486_reg ( .D(n7052), .CK(clk), .RN(n7987), .SN(1'b1), .Q(n12420)
         );
  DFFSRX1 g4489_reg ( .D(n7053), .CK(clk), .RN(n7987), .SN(1'b1), .Q(n12421)
         );
  DFFSRX1 g4492_reg ( .D(n7054), .CK(clk), .RN(n7987), .SN(1'b1), .Q(n12424)
         );
  DFFSRX1 g4504_reg ( .D(n7189), .CK(clk), .RN(n7987), .SN(1'b1), .Q(g4504) );
  DFFSRX1 g4512_reg ( .D(n7064), .CK(clk), .RN(n8078), .SN(1'b1), .Q(n12417)
         );
  DFFSRX1 g4372_reg ( .D(n7190), .CK(clk), .RN(n8078), .SN(1'b1), .Q(n12440), 
        .QN(n7844) );
  DFFSRX1 g4414_reg ( .D(n7185), .CK(clk), .RN(n8078), .SN(1'b1), .Q(g7257), 
        .QN(n5285) );
  DFFSRX1 g1_reg ( .D(n7186), .CK(clk), .RN(n8076), .SN(1'b1), .Q(g12832) );
  DFFSRX1 g4519_reg ( .D(n7188), .CK(clk), .RN(n7988), .SN(1'b1), .Q(g4519) );
  DFFSRX1 g4520_reg ( .D(g4519), .CK(clk), .RN(n7988), .SN(1'b1), .Q(n12416)
         );
  DFFSRX1 g4549_reg ( .D(n7176), .CK(clk), .RN(n8078), .SN(1'b1), .Q(g4549) );
  DFFSRX1 g4552_reg ( .D(n7065), .CK(clk), .RN(n8078), .SN(1'b1), .Q(n12407)
         );
  DFFSRX1 g4570_reg ( .D(n7175), .CK(clk), .RN(n8078), .SN(1'b1), .Q(g4570) );
  DFFSRX1 g4571_reg ( .D(g4570), .CK(clk), .RN(n8078), .SN(1'b1), .Q(n12157)
         );
  DFFSRX1 g4555_reg ( .D(n7083), .CK(clk), .RN(n7985), .SN(1'b1), .Q(n12413)
         );
  DFFSRX1 g4558_reg ( .D(n7055), .CK(clk), .RN(n7985), .SN(1'b1), .Q(n12412)
         );
  DFFSRX1 g4561_reg ( .D(n7056), .CK(clk), .RN(n7985), .SN(1'b1), .Q(n12411)
         );
  DFFSRX1 g2844_reg ( .D(n7138), .CK(clk), .RN(n8080), .SN(1'b1), .Q(n12685), 
        .QN(n7784) );
  DFFSRX1 g554_reg ( .D(n7096), .CK(clk), .RN(n8083), .SN(1'b1), .Q(n12924), 
        .QN(n7816) );
  DFFSRX1 g6711_reg ( .D(n7072), .CK(clk), .RN(n8033), .SN(1'b1), .Q(g17871), 
        .QN(n5253) );
  DFFSRX1 g6715_reg ( .D(g17871), .CK(clk), .RN(n8033), .SN(1'b1), .Q(g14749), 
        .QN(n5270) );
  DFFSRX1 g6494_reg ( .D(n7073), .CK(clk), .RN(n8033), .SN(1'b1), .Q(n12187), 
        .QN(n7771) );
  DFFSRX1 g6444_reg ( .D(n7162), .CK(clk), .RN(n8033), .SN(1'b1), .Q(n12188)
         );
  DFFSRX1 g4894_reg ( .D(n7166), .CK(clk), .RN(n8032), .SN(1'b1), .Q(n12306)
         );
  DFFSRX1 g4888_reg ( .D(n7132), .CK(clk), .RN(n8032), .SN(1'b1), .Q(n12391), 
        .QN(n7700) );
  DFFSRX1 g807_reg ( .D(n6865), .CK(clk), .RN(n8083), .SN(1'b1), .Q(n12925), 
        .QN(n7573) );
  DFFSRX1 g164_reg ( .D(n6864), .CK(clk), .RN(n8083), .SN(1'b1), .Q(n12900), 
        .QN(n7607) );
  DFFSRX1 g168_reg ( .D(n6863), .CK(clk), .RN(n8026), .SN(1'b1), .Q(n12901), 
        .QN(n7634) );
  DFFSRX1 g174_reg ( .D(n6862), .CK(clk), .RN(n8026), .SN(1'b1), .Q(n12902) );
  DFFSRX1 g854_reg ( .D(n6861), .CK(clk), .RN(n8025), .SN(1'b1), .Q(n12489) );
  DFFSRX1 g862_reg ( .D(n6860), .CK(clk), .RN(n8022), .SN(1'b1), .Q(n12769), 
        .QN(n7528) );
  DFFSRX1 g890_reg ( .D(n6859), .CK(clk), .RN(n8022), .SN(1'b1), .Q(n12771), 
        .QN(n7258) );
  DFFSRX1 g896_reg ( .D(n6858), .CK(clk), .RN(n8022), .SN(1'b1), .QN(n12770)
         );
  DFFSRX1 g956_reg ( .D(n6857), .CK(clk), .RN(n8022), .SN(1'b1), .Q(n7362), 
        .QN(n13035) );
  DFFSRX1 g962_reg ( .D(n6856), .CK(clk), .RN(n8021), .SN(1'b1), .Q(n13017), 
        .QN(n7640) );
  DFFSRX1 g969_reg ( .D(n6855), .CK(clk), .RN(n8020), .SN(1'b1), .Q(n13068), 
        .QN(n7609) );
  DFFSRX1 g976_reg ( .D(n6854), .CK(clk), .RN(n8019), .SN(1'b1), .Q(n13042) );
  DFFSRX1 g979_reg ( .D(n6853), .CK(clk), .RN(n8022), .SN(1'b1), .Q(n13074), 
        .QN(n7266) );
  DFFSRX1 g1996_reg ( .D(n6852), .CK(clk), .RN(n8005), .SN(1'b1), .Q(n12819), 
        .QN(n7403) );
  DFFSRX1 g2089_reg ( .D(n6851), .CK(clk), .RN(n8000), .SN(1'b1), .Q(n12810)
         );
  DFFSRX1 g2093_reg ( .D(n6850), .CK(clk), .RN(n7999), .SN(1'b1), .Q(n12798), 
        .QN(n7515) );
  DFFSRX1 g2098_reg ( .D(n6849), .CK(clk), .RN(n7999), .SN(1'b1), .Q(n7601), 
        .QN(n12797) );
  DFFSRX1 g2102_reg ( .D(n6848), .CK(clk), .RN(n7999), .SN(1'b1), .Q(n12796), 
        .QN(n7580) );
  DFFSRX1 g2108_reg ( .D(n6847), .CK(clk), .RN(n7998), .SN(1'b1), .Q(n12795)
         );
  DFFSRX1 g2112_reg ( .D(n6846), .CK(clk), .RN(n7998), .SN(1'b1), .QN(n7240)
         );
  DFFSRX1 g2116_reg ( .D(n6845), .CK(clk), .RN(n7998), .SN(1'b1), .Q(n12794), 
        .QN(n7307) );
  DFFSRX1 g2122_reg ( .D(n6844), .CK(clk), .RN(n7998), .SN(1'b1), .QN(n7651)
         );
  DFFSRX1 g2126_reg ( .D(n6843), .CK(clk), .RN(n7998), .SN(1'b1), .QN(n7215)
         );
  DFFSRX1 g2153_reg ( .D(n6842), .CK(clk), .RN(n7989), .SN(1'b1), .Q(n12792), 
        .QN(n7265) );
  DFFSRX1 g2246_reg ( .D(n6841), .CK(clk), .RN(n7989), .SN(1'b1), .Q(n12788)
         );
  DFFSRX1 g2250_reg ( .D(n6840), .CK(clk), .RN(n8011), .SN(1'b1), .Q(n7432), 
        .QN(n12775) );
  DFFSRX1 g2255_reg ( .D(n6839), .CK(clk), .RN(n8011), .SN(1'b1), .Q(n12774), 
        .QN(n7765) );
  DFFSRX1 g2848_reg ( .D(n6838), .CK(clk), .RN(n8080), .SN(1'b1), .Q(n12683), 
        .QN(n7741) );
  DFFSRX1 g2864_reg ( .D(n6837), .CK(clk), .RN(n7985), .SN(1'b1), .Q(n12671), 
        .QN(n7744) );
  DFFSRX1 g2898_reg ( .D(n6836), .CK(clk), .RN(n8080), .SN(1'b1), .Q(n12665), 
        .QN(n7742) );
  DFFSRX1 g2902_reg ( .D(n6835), .CK(clk), .RN(n8082), .SN(1'b1), .Q(n12660), 
        .QN(n7670) );
  DFFSRX1 g2907_reg ( .D(n6834), .CK(clk), .RN(n8079), .SN(1'b1), .Q(n12658)
         );
  DFFSRX1 g2912_reg ( .D(n6833), .CK(clk), .RN(n8079), .SN(1'b1), .Q(n12656), 
        .QN(n7706) );
  DFFSRX1 g2917_reg ( .D(n6832), .CK(clk), .RN(n8082), .SN(1'b1), .Q(n12655), 
        .QN(n7671) );
  DFFSRX1 g2922_reg ( .D(n6831), .CK(clk), .RN(n8079), .SN(1'b1), .Q(n12654)
         );
  DFFSRX1 g2927_reg ( .D(n6830), .CK(clk), .RN(n8082), .SN(1'b1), .Q(n12652), 
        .QN(n7766) );
  DFFSRX1 g2936_reg ( .D(n6829), .CK(clk), .RN(n8058), .SN(1'b1), .Q(n12651), 
        .QN(n7707) );
  DFFSRX1 g2941_reg ( .D(n6828), .CK(clk), .RN(n8082), .SN(1'b1), .Q(n12647), 
        .QN(n7672) );
  DFFSRX1 g2946_reg ( .D(n6827), .CK(clk), .RN(n8057), .SN(1'b1), .Q(n7598), 
        .QN(n12663) );
  DFFSRX1 g2950_reg ( .D(n6826), .CK(clk), .RN(n8057), .SN(1'b1), .Q(n12646), 
        .QN(n7708) );
  DFFSRX1 g2955_reg ( .D(n6825), .CK(clk), .RN(n8081), .SN(1'b1), .Q(n12645), 
        .QN(n7673) );
  DFFSRX1 g2960_reg ( .D(n6824), .CK(clk), .RN(n8057), .SN(1'b1), .Q(n12644)
         );
  DFFSRX1 g2965_reg ( .D(n6823), .CK(clk), .RN(n8081), .SN(1'b1), .Q(n12643), 
        .QN(n7787) );
  DFFSRX1 g2970_reg ( .D(n6822), .CK(clk), .RN(n8057), .SN(1'b1), .Q(n12659), 
        .QN(n7709) );
  DFFSRX1 g2975_reg ( .D(n6821), .CK(clk), .RN(n8081), .SN(1'b1), .Q(n12642), 
        .QN(n7674) );
  DFFSRX1 g2980_reg ( .D(n6820), .CK(clk), .RN(n8079), .SN(1'b1), .Q(n12641), 
        .QN(n7835) );
  DFFSRX1 g2988_reg ( .D(n6819), .CK(clk), .RN(n8079), .SN(1'b1), .Q(n12668), 
        .QN(n7759) );
  DFFSRX1 g2868_reg ( .D(n6818), .CK(clk), .RN(n7985), .SN(1'b1), .Q(n12669)
         );
  DFFSRX1 g2873_reg ( .D(n6817), .CK(clk), .RN(n7985), .SN(1'b1), .Q(n12667), 
        .QN(n7350) );
  DFFSRX1 g3003_reg ( .D(n6816), .CK(clk), .RN(n8081), .SN(1'b1), .QN(n7827)
         );
  DFFSRX1 g3096_reg ( .D(n6815), .CK(clk), .RN(n8081), .SN(1'b1), .Q(g8277), 
        .QN(n7975) );
  DFFSRX1 g3106_reg ( .D(n6814), .CK(clk), .RN(n8081), .SN(1'b1), .QN(n12602)
         );
  DFFSRX1 g3115_reg ( .D(n6813), .CK(clk), .RN(n8081), .SN(1'b1), .Q(n12674), 
        .QN(n7229) );
  DFFSRX1 g3119_reg ( .D(n6812), .CK(clk), .RN(n8081), .SN(1'b1), .Q(n12598), 
        .QN(n7558) );
  DFFSRX1 g3125_reg ( .D(n6811), .CK(clk), .RN(n8030), .SN(1'b1), .QN(n12597)
         );
  DFFSRX1 g3129_reg ( .D(n6810), .CK(clk), .RN(n8081), .SN(1'b1), .QN(n12689)
         );
  DFFSRX1 g3133_reg ( .D(n6809), .CK(clk), .RN(n8069), .SN(1'b1), .Q(n12596), 
        .QN(n7559) );
  DFFSRX1 g3139_reg ( .D(n6808), .CK(clk), .RN(n8068), .SN(1'b1), .Q(n12595)
         );
  DFFSRX1 g3143_reg ( .D(n6807), .CK(clk), .RN(n8069), .SN(1'b1), .QN(n7644)
         );
  DFFSRX1 g3155_reg ( .D(n6806), .CK(clk), .RN(n8068), .SN(1'b1), .Q(n12592), 
        .QN(n7301) );
  DFFSRX1 g3161_reg ( .D(n6805), .CK(clk), .RN(n8068), .SN(1'b1), .Q(n12591), 
        .QN(n7564) );
  DFFSRX1 g3167_reg ( .D(n6804), .CK(clk), .RN(n8068), .SN(1'b1), .Q(n12600), 
        .QN(n7217) );
  DFFSRX1 g3171_reg ( .D(n6803), .CK(clk), .RN(n8068), .SN(1'b1), .Q(n12601)
         );
  DFFSRX1 g3179_reg ( .D(n6802), .CK(clk), .RN(n8068), .SN(1'b1), .Q(n12636), 
        .QN(n7480) );
  DFFSRX1 g3092_reg ( .D(n6801), .CK(clk), .RN(n8081), .SN(1'b1), .Q(g8215), 
        .QN(n489) );
  DFFSRX1 g3187_reg ( .D(n6800), .CK(clk), .RN(n8055), .SN(1'b1), .Q(n12616)
         );
  DFFSRX1 g3215_reg ( .D(n6799), .CK(clk), .RN(n8055), .SN(1'b1), .Q(n12615)
         );
  DFFSRX1 g3231_reg ( .D(n6798), .CK(clk), .RN(n8068), .SN(1'b1), .Q(n12613)
         );
  DFFSRX1 g3247_reg ( .D(n6797), .CK(clk), .RN(n8056), .SN(1'b1), .Q(n7225) );
  DFFSRX1 g3251_reg ( .D(n6796), .CK(clk), .RN(n8056), .SN(1'b1), .Q(n12626)
         );
  DFFSRX1 g3255_reg ( .D(n6795), .CK(clk), .RN(n8056), .SN(1'b1), .Q(n12620)
         );
  DFFSRX1 g3259_reg ( .D(n6794), .CK(clk), .RN(n8056), .SN(1'b1), .Q(n12621), 
        .QN(n7788) );
  DFFSRX1 g3263_reg ( .D(n6793), .CK(clk), .RN(n8049), .SN(1'b1), .Q(n12614)
         );
  DFFSRX1 g3333_reg ( .D(n6792), .CK(clk), .RN(n8068), .SN(1'b1), .Q(n12587), 
        .QN(n7781) );
  DFFSRX1 g3338_reg ( .D(n6791), .CK(clk), .RN(n8067), .SN(1'b1), .Q(n12635), 
        .QN(n7422) );
  DFFSRX1 g3343_reg ( .D(n6790), .CK(clk), .RN(n8067), .SN(1'b1), .QN(n7652)
         );
  DFFSRX1 g3347_reg ( .D(n6789), .CK(clk), .RN(n8067), .SN(1'b1), .Q(n12586), 
        .QN(n7624) );
  DFFSRX1 g4939_reg ( .D(n6788), .CK(clk), .RN(n8067), .SN(1'b1), .Q(n12302), 
        .QN(n7779) );
  DFFSRX1 g4966_reg ( .D(n6787), .CK(clk), .RN(n8037), .SN(1'b1), .Q(n7363), 
        .QN(n12610) );
  DFFSRX1 g4975_reg ( .D(n6786), .CK(clk), .RN(n8037), .SN(1'b1), .Q(n7247), 
        .QN(n12612) );
  DFFSRX1 g4899_reg ( .D(n6785), .CK(clk), .RN(n8032), .SN(1'b1), .Q(n7379), 
        .QN(n12611) );
  DFFSRX1 g4907_reg ( .D(n6784), .CK(clk), .RN(n8032), .SN(1'b1), .Q(n12390)
         );
  DFFSRX1 g4912_reg ( .D(n6783), .CK(clk), .RN(n8031), .SN(1'b1), .Q(n12389)
         );
  DFFSRX1 g4927_reg ( .D(n6782), .CK(clk), .RN(n8031), .SN(1'b1), .Q(n12388), 
        .QN(n7746) );
  DFFSRX1 g4933_reg ( .D(n6781), .CK(clk), .RN(n8030), .SN(1'b1), .Q(n7499), 
        .QN(n12604) );
  DFFSRX1 g4581_reg ( .D(n6780), .CK(clk), .RN(n8075), .SN(1'b1), .Q(n12425), 
        .QN(n7685) );
  DFFSRX1 g4584_reg ( .D(n6779), .CK(clk), .RN(n8075), .SN(1'b1), .Q(n7359), 
        .QN(n12446) );
  DFFSRX1 g4593_reg ( .D(n6778), .CK(clk), .RN(n8075), .SN(1'b1), .Q(n7355), 
        .QN(n12442) );
  DFFSRX1 g4601_reg ( .D(n6777), .CK(clk), .RN(n8075), .SN(1'b1), .Q(n7410), 
        .QN(n12443) );
  DFFSRX1 g4608_reg ( .D(n6776), .CK(clk), .RN(n8075), .SN(1'b1), .QN(n12445)
         );
  DFFSRX1 g4616_reg ( .D(n6775), .CK(clk), .RN(n8075), .SN(1'b1), .QN(n12444)
         );
  DFFSRX1 g4621_reg ( .D(n6774), .CK(clk), .RN(n8075), .SN(1'b1), .Q(n7413), 
        .QN(n12455) );
  DFFSRX1 g4628_reg ( .D(n6773), .CK(clk), .RN(n8028), .SN(1'b1), .Q(n7277), 
        .QN(n12454) );
  DFFSRX1 g4633_reg ( .D(n6772), .CK(clk), .RN(n8028), .SN(1'b1), .Q(n7276), 
        .QN(n12385) );
  DFFSRX1 g4643_reg ( .D(n6771), .CK(clk), .RN(n8075), .SN(1'b1), .Q(n7245), 
        .QN(n12450) );
  DFFSRX1 g4639_reg ( .D(n6770), .CK(clk), .RN(n8028), .SN(1'b1), .QN(n12456)
         );
  DFFSRX1 g4646_reg ( .D(n6769), .CK(clk), .RN(n8075), .SN(1'b1), .Q(n12995), 
        .QN(n7608) );
  DFFSRX1 g4653_reg ( .D(n6768), .CK(clk), .RN(n8074), .SN(1'b1), .Q(n12999), 
        .QN(n7577) );
  DFFSRX1 g4659_reg ( .D(n6767), .CK(clk), .RN(n8074), .SN(1'b1), .Q(n7433), 
        .QN(n12996) );
  DFFSRX1 g4664_reg ( .D(n6766), .CK(clk), .RN(n8074), .SN(1'b1), .QN(n7653)
         );
  DFFSRX1 g4669_reg ( .D(n6765), .CK(clk), .RN(n8074), .SN(1'b1), .Q(n12998), 
        .QN(n7546) );
  DFFSRX1 g4674_reg ( .D(n6764), .CK(clk), .RN(n8075), .SN(1'b1), .Q(n6763), 
        .QN(n12404) );
  DFFSRX1 g4681_reg ( .D(n6763), .CK(clk), .RN(n8075), .SN(1'b1), .Q(n4749), 
        .QN(n12403) );
  DFFSRX1 g4688_reg ( .D(n4749), .CK(clk), .RN(n8075), .SN(1'b1), .Q(n7360), 
        .QN(n12405) );
  DFFSRX1 g5462_reg ( .D(n6762), .CK(clk), .RN(n8043), .SN(1'b1), .Q(n7578), 
        .QN(n12239) );
  DFFSRX1 g5471_reg ( .D(n6761), .CK(clk), .RN(n8043), .SN(1'b1), .Q(n12678), 
        .QN(n7230) );
  DFFSRX1 g5475_reg ( .D(n6760), .CK(clk), .RN(n8043), .SN(1'b1), .Q(n12234), 
        .QN(n7560) );
  DFFSRX1 g5481_reg ( .D(n6759), .CK(clk), .RN(n8039), .SN(1'b1), .QN(n12233)
         );
  DFFSRX1 g5485_reg ( .D(n6758), .CK(clk), .RN(n8043), .SN(1'b1), .Q(n7599), 
        .QN(n12696) );
  DFFSRX1 g5489_reg ( .D(n6757), .CK(clk), .RN(n8043), .SN(1'b1), .Q(n12232), 
        .QN(n7561) );
  DFFSRX1 g5495_reg ( .D(n6756), .CK(clk), .RN(n8042), .SN(1'b1), .Q(n12231)
         );
  DFFSRX1 g5499_reg ( .D(n6755), .CK(clk), .RN(n8043), .SN(1'b1), .Q(n12695), 
        .QN(n7622) );
  DFFSRX1 g5511_reg ( .D(n6754), .CK(clk), .RN(n8043), .SN(1'b1), .QN(n12230)
         );
  DFFSRX1 g5517_reg ( .D(n6753), .CK(clk), .RN(n8043), .SN(1'b1), .Q(n7425), 
        .QN(n12229) );
  DFFSRX1 g5523_reg ( .D(n6752), .CK(clk), .RN(n8043), .SN(1'b1), .Q(n12236), 
        .QN(n7259) );
  DFFSRX1 g5527_reg ( .D(n6751), .CK(clk), .RN(n8043), .SN(1'b1), .QN(n12237)
         );
  DFFSRX1 g5535_reg ( .D(n6750), .CK(clk), .RN(n8043), .SN(1'b1), .Q(n12240), 
        .QN(n7481) );
  DFFSRX1 g5567_reg ( .D(n6749), .CK(clk), .RN(n8042), .SN(1'b1), .Q(n12368)
         );
  DFFSRX1 g5571_reg ( .D(n6748), .CK(clk), .RN(n8042), .SN(1'b1), .Q(n12355)
         );
  DFFSRX1 g5587_reg ( .D(n6747), .CK(clk), .RN(n8042), .SN(1'b1), .Q(n12354)
         );
  DFFSRX1 g5603_reg ( .D(n6746), .CK(clk), .RN(n8042), .SN(1'b1), .Q(n7226) );
  DFFSRX1 g5607_reg ( .D(n6745), .CK(clk), .RN(n8041), .SN(1'b1), .Q(n12365)
         );
  DFFSRX1 g5611_reg ( .D(n6744), .CK(clk), .RN(n8041), .SN(1'b1), .Q(n12358)
         );
  DFFSRX1 g5615_reg ( .D(n6743), .CK(clk), .RN(n8041), .SN(1'b1), .Q(n12360), 
        .QN(n7790) );
  DFFSRX1 g5619_reg ( .D(n6742), .CK(clk), .RN(n8041), .SN(1'b1), .Q(n12371)
         );
  DFFSRX1 g5623_reg ( .D(n6741), .CK(clk), .RN(n8041), .SN(1'b1), .Q(g17580), 
        .QN(n5778) );
  DFFSRX1 g5630_reg ( .D(g17580), .CK(clk), .RN(n8041), .SN(1'b1), .Q(g17604), 
        .QN(n7817) );
  DFFSRX1 g5659_reg ( .D(n6740), .CK(clk), .RN(n8039), .SN(1'b1), .Q(g12300)
         );
  DFFSRX1 g5637_reg ( .D(n6739), .CK(clk), .RN(n8039), .SN(1'b1), .Q(g14694)
         );
  DFFSRX1 g5666_reg ( .D(n6738), .CK(clk), .RN(n8039), .SN(1'b1), .Q(g17711), 
        .QN(n5779) );
  DFFSRX1 g5681_reg ( .D(g14635), .CK(clk), .RN(n8039), .SN(1'b1), .Q(g17678)
         );
  DFFSRX1 g5685_reg ( .D(g17678), .CK(clk), .RN(n8039), .SN(1'b1), .Q(n12367), 
        .QN(n7791) );
  DFFSRX1 g5689_reg ( .D(n6736), .CK(clk), .RN(n8040), .SN(1'b1), .Q(n7415), 
        .QN(n12356) );
  DFFSRX1 g5694_reg ( .D(n6735), .CK(clk), .RN(n8040), .SN(1'b1), .QN(n7658)
         );
  DFFSRX1 g5698_reg ( .D(n6734), .CK(clk), .RN(n8040), .SN(1'b1), .Q(n12380), 
        .QN(n7627) );
  DFFSRX1 g5703_reg ( .D(n6733), .CK(clk), .RN(n8040), .SN(1'b1), .Q(n7295), 
        .QN(n12382) );
  DFFSRX1 g5644_reg ( .D(n6732), .CK(clk), .RN(n8039), .SN(1'b1), .Q(n12381), 
        .QN(n7545) );
  DFFSRX1 g5654_reg ( .D(n6731), .CK(clk), .RN(n8039), .SN(1'b1), .Q(g13049)
         );
  DFFSRX1 g4826_reg ( .D(n6730), .CK(clk), .RN(n8038), .SN(1'b1), .Q(n7504), 
        .QN(n12395) );
  DFFSRX1 g4836_reg ( .D(n6729), .CK(clk), .RN(n8069), .SN(1'b1), .Q(n7431), 
        .QN(n12392) );
  DFFSRX1 g4843_reg ( .D(n6728), .CK(clk), .RN(n8069), .SN(1'b1), .Q(n12607), 
        .QN(n7576) );
  DFFSRX1 g4849_reg ( .D(n6727), .CK(clk), .RN(n8069), .SN(1'b1), .Q(n7434), 
        .QN(n12605) );
  DFFSRX1 g4983_reg ( .D(n6726), .CK(clk), .RN(n8037), .SN(1'b1), .Q(n7250), 
        .QN(n12609) );
  DFFSRX1 g4991_reg ( .D(n6725), .CK(clk), .RN(n8037), .SN(1'b1), .Q(n7411), 
        .QN(n12608) );
  DFFSRX1 g4854_reg ( .D(n6724), .CK(clk), .RN(n8069), .SN(1'b1), .QN(n7654)
         );
  DFFSRX1 g4859_reg ( .D(n6723), .CK(clk), .RN(n8069), .SN(1'b1), .Q(n12606), 
        .QN(n7541) );
  DFFSRX1 g4864_reg ( .D(n6722), .CK(clk), .RN(n8069), .SN(1'b1), .Q(n4770), 
        .QN(n12603) );
  DFFSRX1 g4871_reg ( .D(n4770), .CK(clk), .RN(n8069), .SN(1'b1), .Q(n4771), 
        .QN(n12549) );
  DFFSRX1 g4878_reg ( .D(n4771), .CK(clk), .RN(n8069), .SN(1'b1), .Q(n12524), 
        .QN(n7285) );
  DFFSRX1 g3352_reg ( .D(n6721), .CK(clk), .RN(n8067), .SN(1'b1), .Q(n12632), 
        .QN(n7242) );
  DFFSRX1 g3288_reg ( .D(n6720), .CK(clk), .RN(n8048), .SN(1'b1), .Q(n12633), 
        .QN(n7361) );
  DFFSRX1 g3298_reg ( .D(n6719), .CK(clk), .RN(n8048), .SN(1'b1), .Q(g14421)
         );
  DFFSRX1 g3303_reg ( .D(n6718), .CK(clk), .RN(n8048), .SN(1'b1), .Q(g11349)
         );
  DFFSRX1 g3310_reg ( .D(n6717), .CK(clk), .RN(n8048), .SN(1'b1), .Q(g16718), 
        .QN(n5824) );
  DFFSRX1 g3267_reg ( .D(n6716), .CK(clk), .RN(n8048), .SN(1'b1), .Q(g16603), 
        .QN(n5825) );
  DFFSRX1 g3274_reg ( .D(g16603), .CK(clk), .RN(n8048), .SN(1'b1), .Q(g16624), 
        .QN(n7837) );
  DFFSRX1 g3281_reg ( .D(n6715), .CK(clk), .RN(n8048), .SN(1'b1), .Q(g13895), 
        .QN(n5826) );
  DFFSRX1 g3325_reg ( .D(g13865), .CK(clk), .RN(n8048), .SN(1'b1), .Q(g16686)
         );
  DFFSRX1 g3329_reg ( .D(g16686), .CK(clk), .RN(n8048), .SN(1'b1), .Q(n12630)
         );
  DFFSRX1 g3447_reg ( .D(n6713), .CK(clk), .RN(n8065), .SN(1'b1), .Q(g8342), 
        .QN(n7973) );
  DFFSRX1 g3457_reg ( .D(n6712), .CK(clk), .RN(n8064), .SN(1'b1), .Q(n12572), 
        .QN(n7526) );
  DFFSRX1 g3466_reg ( .D(n6711), .CK(clk), .RN(n8067), .SN(1'b1), .Q(n12673), 
        .QN(n7322) );
  DFFSRX1 g3470_reg ( .D(n6710), .CK(clk), .RN(n8067), .SN(1'b1), .QN(n7398)
         );
  DFFSRX1 g3476_reg ( .D(n6709), .CK(clk), .RN(n8067), .SN(1'b1), .Q(n12544)
         );
  DFFSRX1 g3480_reg ( .D(n6708), .CK(clk), .RN(n8067), .SN(1'b1), .QN(n7643)
         );
  DFFSRX1 g3484_reg ( .D(n6707), .CK(clk), .RN(n8067), .SN(1'b1), .Q(n12543), 
        .QN(n7581) );
  DFFSRX1 g3490_reg ( .D(n6706), .CK(clk), .RN(n8066), .SN(1'b1), .Q(n12542)
         );
  DFFSRX1 g3494_reg ( .D(n6705), .CK(clk), .RN(n8067), .SN(1'b1), .QN(n7333)
         );
  DFFSRX1 g3506_reg ( .D(n6704), .CK(clk), .RN(n8066), .SN(1'b1), .Q(n12535), 
        .QN(n7298) );
  DFFSRX1 g3512_reg ( .D(n6703), .CK(clk), .RN(n8066), .SN(1'b1), .Q(n12534), 
        .QN(n7565) );
  DFFSRX1 g3518_reg ( .D(n6702), .CK(clk), .RN(n8066), .SN(1'b1), .Q(n12546), 
        .QN(n7220) );
  DFFSRX1 g3522_reg ( .D(n6701), .CK(clk), .RN(n8066), .SN(1'b1), .Q(n12547), 
        .QN(n7267) );
  DFFSRX1 g3530_reg ( .D(n6700), .CK(clk), .RN(n8066), .SN(1'b1), .Q(n12574), 
        .QN(n7507) );
  DFFSRX1 g3443_reg ( .D(n6699), .CK(clk), .RN(n8065), .SN(1'b1), .Q(g8279), 
        .QN(n524) );
  DFFSRX1 g3562_reg ( .D(n6698), .CK(clk), .RN(n8049), .SN(1'b1), .Q(n12567)
         );
  DFFSRX1 g3566_reg ( .D(n6697), .CK(clk), .RN(n8049), .SN(1'b1), .Q(n12556)
         );
  DFFSRX1 g3582_reg ( .D(n6696), .CK(clk), .RN(n8049), .SN(1'b1), .Q(n12555)
         );
  DFFSRX1 g3598_reg ( .D(n6695), .CK(clk), .RN(n8049), .SN(1'b1), .Q(n7279) );
  DFFSRX1 g3602_reg ( .D(n6694), .CK(clk), .RN(n8050), .SN(1'b1), .Q(n12564)
         );
  DFFSRX1 g3606_reg ( .D(n6693), .CK(clk), .RN(n8050), .SN(1'b1), .Q(n12558)
         );
  DFFSRX1 g3610_reg ( .D(n6692), .CK(clk), .RN(n8066), .SN(1'b1), .Q(n12561), 
        .QN(n7792) );
  DFFSRX1 g3614_reg ( .D(n6691), .CK(clk), .RN(n8066), .SN(1'b1), .Q(n12554)
         );
  DFFSRX1 g3689_reg ( .D(n6690), .CK(clk), .RN(n8065), .SN(1'b1), .Q(n12573), 
        .QN(n7374) );
  DFFSRX1 g3694_reg ( .D(n6689), .CK(clk), .RN(n8065), .SN(1'b1), .QN(n12529)
         );
  DFFSRX1 g3698_reg ( .D(n6688), .CK(clk), .RN(n8064), .SN(1'b1), .Q(n12530)
         );
  DFFSRX1 g3703_reg ( .D(n6687), .CK(clk), .RN(n8064), .SN(1'b1), .Q(n12571), 
        .QN(n7274) );
  DFFSRX1 g3798_reg ( .D(n6686), .CK(clk), .RN(n8063), .SN(1'b1), .Q(g8398), 
        .QN(n3810) );
  DFFSRX1 g3808_reg ( .D(n6685), .CK(clk), .RN(n8063), .SN(1'b1), .Q(n12501), 
        .QN(n7513) );
  DFFSRX1 g3817_reg ( .D(n6684), .CK(clk), .RN(n8063), .SN(1'b1), .Q(n12672), 
        .QN(n7620) );
  DFFSRX1 g3821_reg ( .D(n6683), .CK(clk), .RN(n8063), .SN(1'b1), .Q(n12496), 
        .QN(n7562) );
  DFFSRX1 g3827_reg ( .D(n6682), .CK(clk), .RN(n8030), .SN(1'b1), .QN(n7655)
         );
  DFFSRX1 g3831_reg ( .D(n6681), .CK(clk), .RN(n8063), .SN(1'b1), .QN(n7645)
         );
  DFFSRX1 g3835_reg ( .D(n6680), .CK(clk), .RN(n8063), .SN(1'b1), .Q(n12495), 
        .QN(n7563) );
  DFFSRX1 g3841_reg ( .D(n6679), .CK(clk), .RN(n8062), .SN(1'b1), .Q(n12494)
         );
  DFFSRX1 g3845_reg ( .D(n6678), .CK(clk), .RN(n8063), .SN(1'b1), .QN(n7334)
         );
  DFFSRX1 g3857_reg ( .D(n6677), .CK(clk), .RN(n8063), .SN(1'b1), .Q(n12493), 
        .QN(n7299) );
  DFFSRX1 g3863_reg ( .D(n6676), .CK(clk), .RN(n8063), .SN(1'b1), .Q(n12492), 
        .QN(n7566) );
  DFFSRX1 g3869_reg ( .D(n6675), .CK(clk), .RN(n8062), .SN(1'b1), .Q(n12498), 
        .QN(n7221) );
  DFFSRX1 g3873_reg ( .D(n6674), .CK(clk), .RN(n8062), .SN(1'b1), .Q(n12499), 
        .QN(n7268) );
  DFFSRX1 g3881_reg ( .D(n6673), .CK(clk), .RN(n8062), .SN(1'b1), .Q(n12526), 
        .QN(n7508) );
  DFFSRX1 g3794_reg ( .D(n6672), .CK(clk), .RN(n8064), .SN(1'b1), .Q(g8344), 
        .QN(n7984) );
  DFFSRX1 g3913_reg ( .D(n6671), .CK(clk), .RN(n8051), .SN(1'b1), .Q(n12518)
         );
  DFFSRX1 g3917_reg ( .D(n6670), .CK(clk), .RN(n8051), .SN(1'b1), .Q(n12507)
         );
  DFFSRX1 g3933_reg ( .D(n6669), .CK(clk), .RN(n8050), .SN(1'b1), .Q(n12506)
         );
  DFFSRX1 g3949_reg ( .D(n6668), .CK(clk), .RN(n8050), .SN(1'b1), .Q(n7280) );
  DFFSRX1 g3953_reg ( .D(n6667), .CK(clk), .RN(n8051), .SN(1'b1), .Q(n12515)
         );
  DFFSRX1 g3957_reg ( .D(n6666), .CK(clk), .RN(n8051), .SN(1'b1), .Q(n12509)
         );
  DFFSRX1 g3961_reg ( .D(n6665), .CK(clk), .RN(n8051), .SN(1'b1), .Q(n12512), 
        .QN(n7793) );
  DFFSRX1 g3965_reg ( .D(n6664), .CK(clk), .RN(n8049), .SN(1'b1), .Q(n12505)
         );
  DFFSRX1 g4035_reg ( .D(n6663), .CK(clk), .RN(n8062), .SN(1'b1), .Q(n12486), 
        .QN(n7782) );
  DFFSRX1 g4040_reg ( .D(n6662), .CK(clk), .RN(n8062), .SN(1'b1), .Q(n12525), 
        .QN(n7369) );
  DFFSRX1 g4045_reg ( .D(n6661), .CK(clk), .RN(n8062), .SN(1'b1), .QN(n12484)
         );
  DFFSRX1 g4049_reg ( .D(n6660), .CK(clk), .RN(n8062), .SN(1'b1), .Q(n12485)
         );
  DFFSRX1 g4054_reg ( .D(n6659), .CK(clk), .RN(n8062), .SN(1'b1), .Q(n12520)
         );
  DFFSRX1 g4057_reg ( .D(n6658), .CK(clk), .RN(n8061), .SN(1'b1), .Q(n12582), 
        .QN(n7384) );
  DFFSRX1 g4122_reg ( .D(n6657), .CK(clk), .RN(n8061), .SN(1'b1), .Q(n12474)
         );
  DFFSRX1 g4141_reg ( .D(n6656), .CK(clk), .RN(n8061), .SN(1'b1), .Q(n12577), 
        .QN(n7676) );
  DFFSRX1 g4082_reg ( .D(n6655), .CK(clk), .RN(n8061), .SN(1'b1), .Q(n12576), 
        .QN(n7340) );
  DFFSRX1 g4087_reg ( .D(n6654), .CK(clk), .RN(n8061), .SN(1'b1), .Q(n12578)
         );
  DFFSRX1 g4093_reg ( .D(n6653), .CK(clk), .RN(n8061), .SN(1'b1), .QN(n7236)
         );
  DFFSRX1 g4098_reg ( .D(n6652), .CK(clk), .RN(n8060), .SN(1'b1), .Q(n12579)
         );
  DFFSRX1 g4072_reg ( .D(n6651), .CK(clk), .RN(n8061), .SN(1'b1), .Q(n12648), 
        .QN(n7231) );
  DFFSRX1 g4064_reg ( .D(n6650), .CK(clk), .RN(n8061), .SN(1'b1), .Q(n12575), 
        .QN(n7269) );
  DFFSRX1 g4076_reg ( .D(n6649), .CK(clk), .RN(n8061), .SN(1'b1), .Q(n12581), 
        .QN(n7330) );
  DFFSRX1 g4104_reg ( .D(n6648), .CK(clk), .RN(n8060), .SN(1'b1), .Q(n12482)
         );
  DFFSRX1 g4108_reg ( .D(n6647), .CK(clk), .RN(n8060), .SN(1'b1), .Q(n12483), 
        .QN(n7839) );
  DFFSRX1 g4145_reg ( .D(n6646), .CK(clk), .RN(n8060), .SN(1'b1), .Q(n12481), 
        .QN(n7341) );
  DFFSRX1 g4112_reg ( .D(n6645), .CK(clk), .RN(n8061), .SN(1'b1), .Q(n7506), 
        .QN(n12580) );
  DFFSRX1 g4116_reg ( .D(n6644), .CK(clk), .RN(n8061), .SN(1'b1), .Q(n12480), 
        .QN(n7840) );
  DFFSRX1 g4119_reg ( .D(n6643), .CK(clk), .RN(n8061), .SN(1'b1), .Q(n12479), 
        .QN(n7838) );
  DFFSRX1 g4153_reg ( .D(n6642), .CK(clk), .RN(n8060), .SN(1'b1), .Q(n12649), 
        .QN(n7339) );
  DFFSRX1 g4164_reg ( .D(n6641), .CK(clk), .RN(n8060), .SN(1'b1), .QN(n7819)
         );
  DFFSRX1 g4172_reg ( .D(n6640), .CK(clk), .RN(n8060), .SN(1'b1), .Q(n12470)
         );
  DFFSRX1 g4176_reg ( .D(n6639), .CK(clk), .RN(n8060), .SN(1'b1), .Q(n12472)
         );
  DFFSRX1 g4146_reg ( .D(n6638), .CK(clk), .RN(n8060), .SN(1'b1), .Q(n12473), 
        .QN(n7712) );
  DFFSRX1 g4180_reg ( .D(n6637), .CK(clk), .RN(n8060), .SN(1'b1), .Q(n12594), 
        .QN(n7516) );
  DFFSRX1 g4197_reg ( .D(g8784), .CK(clk), .RN(n8059), .SN(1'b1), .Q(g8785), 
        .QN(n7863) );
  DFFSRX1 g4204_reg ( .D(g8786), .CK(clk), .RN(n8059), .SN(1'b1), .Q(g8787), 
        .QN(n7864) );
  DFFSRX1 g4207_reg ( .D(g8787), .CK(clk), .RN(n8059), .SN(1'b1), .Q(g8788), 
        .QN(n7861) );
  DFFSRX1 g4210_reg ( .D(g8788), .CK(clk), .RN(n8059), .SN(1'b1), .Q(g8789), 
        .QN(n7862) );
  DFFSRX1 g4213_reg ( .D(n6636), .CK(clk), .RN(n8059), .SN(1'b1), .Q(g8915), 
        .QN(n7824) );
  DFFSRX1 g4216_reg ( .D(g8915), .CK(clk), .RN(n8059), .SN(1'b1), .Q(g8916), 
        .QN(n7825) );
  DFFSRX1 g4222_reg ( .D(g8917), .CK(clk), .RN(n8059), .SN(1'b1), .Q(g8870), 
        .QN(n603) );
  DFFSRX1 g4235_reg ( .D(g8920), .CK(clk), .RN(n8058), .SN(1'b1), .Q(n7455), 
        .QN(n12468) );
  DFFSRX1 g4239_reg ( .D(n6635), .CK(clk), .RN(n8037), .SN(1'b1), .Q(n12466), 
        .QN(n7749) );
  DFFSRX1 g4242_reg ( .D(n6634), .CK(clk), .RN(n8058), .SN(1'b1), .Q(n12463), 
        .QN(n7831) );
  DFFSRX1 g4253_reg ( .D(n6633), .CK(clk), .RN(n8058), .SN(1'b1), .Q(n12469)
         );
  DFFSRX1 g4185_reg ( .D(n6632), .CK(clk), .RN(n8037), .SN(1'b1), .Q(g11770), 
        .QN(n7826) );
  DFFSRX1 g4264_reg ( .D(n6631), .CK(clk), .RN(n8057), .SN(1'b1), .Q(n12461), 
        .QN(n7795) );
  DFFSRX1 g4269_reg ( .D(n6630), .CK(clk), .RN(n8057), .SN(1'b1), .Q(n12459), 
        .QN(n7677) );
  DFFSRX1 g4273_reg ( .D(n6629), .CK(clk), .RN(n8057), .SN(1'b1), .Q(n12467), 
        .QN(n7697) );
  DFFSRX1 g4281_reg ( .D(g8839), .CK(clk), .RN(n8057), .SN(1'b1), .QN(n7650)
         );
  DFFSRX1 g3195_reg ( .D(n6628), .CK(clk), .RN(n8055), .SN(1'b1), .Q(n12617)
         );
  DFFSRX1 g3191_reg ( .D(n6627), .CK(clk), .RN(n8055), .SN(1'b1), .Q(n7278) );
  DFFSRX1 g3203_reg ( .D(n6626), .CK(clk), .RN(n8055), .SN(1'b1), .Q(n12619)
         );
  DFFSRX1 g3199_reg ( .D(n6625), .CK(clk), .RN(n8055), .SN(1'b1), .Q(n12629)
         );
  DFFSRX1 g3211_reg ( .D(n6624), .CK(clk), .RN(n8055), .SN(1'b1), .Q(n12631)
         );
  DFFSRX1 g3207_reg ( .D(n6623), .CK(clk), .RN(n8055), .SN(1'b1), .Q(n12624)
         );
  DFFSRX1 g3219_reg ( .D(n6622), .CK(clk), .RN(n8055), .SN(1'b1), .Q(n12627)
         );
  DFFSRX1 g3223_reg ( .D(n6621), .CK(clk), .RN(n8055), .SN(1'b1), .Q(n12618)
         );
  DFFSRX1 g3227_reg ( .D(n6620), .CK(clk), .RN(n8055), .SN(1'b1), .Q(n12623)
         );
  DFFSRX1 g3235_reg ( .D(n6619), .CK(clk), .RN(n8068), .SN(1'b1), .Q(n12625)
         );
  DFFSRX1 g3239_reg ( .D(n6618), .CK(clk), .RN(n8068), .SN(1'b1), .Q(n12628)
         );
  DFFSRX1 g3243_reg ( .D(n6617), .CK(clk), .RN(n8068), .SN(1'b1), .Q(n12622)
         );
  DFFSRX1 g3538_reg ( .D(n6616), .CK(clk), .RN(n8056), .SN(1'b1), .Q(n12551)
         );
  DFFSRX1 g3546_reg ( .D(n6615), .CK(clk), .RN(n8049), .SN(1'b1), .Q(n12552)
         );
  DFFSRX1 g3542_reg ( .D(n6614), .CK(clk), .RN(n8049), .SN(1'b1), .Q(n7438), 
        .QN(n12553) );
  DFFSRX1 g3554_reg ( .D(n6613), .CK(clk), .RN(n8050), .SN(1'b1), .Q(n12557)
         );
  DFFSRX1 g3550_reg ( .D(n6612), .CK(clk), .RN(n8049), .SN(1'b1), .Q(n12565)
         );
  DFFSRX1 g3558_reg ( .D(n6611), .CK(clk), .RN(n8050), .SN(1'b1), .Q(n7386) );
  DFFSRX1 g3570_reg ( .D(n6610), .CK(clk), .RN(n8049), .SN(1'b1), .Q(n12562)
         );
  DFFSRX1 g3574_reg ( .D(n6609), .CK(clk), .RN(n8049), .SN(1'b1), .Q(n12568)
         );
  DFFSRX1 g3578_reg ( .D(n6608), .CK(clk), .RN(n8049), .SN(1'b1), .Q(n12560)
         );
  DFFSRX1 g3586_reg ( .D(n6607), .CK(clk), .RN(n8066), .SN(1'b1), .Q(n12563)
         );
  DFFSRX1 g3590_reg ( .D(n6606), .CK(clk), .RN(n8066), .SN(1'b1), .Q(n12569)
         );
  DFFSRX1 g3594_reg ( .D(n6605), .CK(clk), .RN(n8066), .SN(1'b1), .Q(n12559)
         );
  DFFSRX1 g3889_reg ( .D(n6604), .CK(clk), .RN(n8056), .SN(1'b1), .Q(n12502)
         );
  DFFSRX1 g3897_reg ( .D(n6603), .CK(clk), .RN(n8050), .SN(1'b1), .Q(n12503)
         );
  DFFSRX1 g3893_reg ( .D(n6602), .CK(clk), .RN(n8050), .SN(1'b1), .Q(n7439), 
        .QN(n12504) );
  DFFSRX1 g3905_reg ( .D(n6601), .CK(clk), .RN(n8051), .SN(1'b1), .Q(n12508)
         );
  DFFSRX1 g3901_reg ( .D(n6600), .CK(clk), .RN(n8050), .SN(1'b1), .Q(n12516)
         );
  DFFSRX1 g3909_reg ( .D(n6599), .CK(clk), .RN(n8051), .SN(1'b1), .Q(n7387) );
  DFFSRX1 g3921_reg ( .D(n6598), .CK(clk), .RN(n8050), .SN(1'b1), .Q(n12513)
         );
  DFFSRX1 g3925_reg ( .D(n6597), .CK(clk), .RN(n8050), .SN(1'b1), .Q(n12519)
         );
  DFFSRX1 g3929_reg ( .D(n6596), .CK(clk), .RN(n8050), .SN(1'b1), .Q(n12511)
         );
  DFFSRX1 g3937_reg ( .D(n6595), .CK(clk), .RN(n8062), .SN(1'b1), .Q(n12514)
         );
  DFFSRX1 g3941_reg ( .D(n6594), .CK(clk), .RN(n8062), .SN(1'b1), .Q(n12522)
         );
  DFFSRX1 g3945_reg ( .D(n6593), .CK(clk), .RN(n8062), .SN(1'b1), .Q(n12510)
         );
  DFFSRX1 g5543_reg ( .D(n6592), .CK(clk), .RN(n8042), .SN(1'b1), .Q(n12352)
         );
  DFFSRX1 g5551_reg ( .D(n6591), .CK(clk), .RN(n8042), .SN(1'b1), .Q(n12353)
         );
  DFFSRX1 g5547_reg ( .D(n6590), .CK(clk), .RN(n8042), .SN(1'b1), .Q(n7440), 
        .QN(n12351) );
  DFFSRX1 g5559_reg ( .D(n6589), .CK(clk), .RN(n8041), .SN(1'b1), .Q(n12357)
         );
  DFFSRX1 g5555_reg ( .D(n6588), .CK(clk), .RN(n8041), .SN(1'b1), .Q(n12366)
         );
  DFFSRX1 g5563_reg ( .D(n6587), .CK(clk), .RN(n8042), .SN(1'b1), .Q(n12362)
         );
  DFFSRX1 g5575_reg ( .D(n6586), .CK(clk), .RN(n8041), .SN(1'b1), .Q(n12364)
         );
  DFFSRX1 g5579_reg ( .D(n6585), .CK(clk), .RN(n8041), .SN(1'b1), .Q(n12370)
         );
  DFFSRX1 g5583_reg ( .D(n6584), .CK(clk), .RN(n8042), .SN(1'b1), .Q(n12359)
         );
  DFFSRX1 g5591_reg ( .D(n6583), .CK(clk), .RN(n8041), .SN(1'b1), .Q(n12363)
         );
  DFFSRX1 g5595_reg ( .D(n6582), .CK(clk), .RN(n8041), .SN(1'b1), .Q(n12369)
         );
  DFFSRX1 g5599_reg ( .D(n6581), .CK(clk), .RN(n8042), .SN(1'b1), .Q(n12361)
         );
  DFFSRX1 g4291_reg ( .D(g9019), .CK(clk), .RN(n8057), .SN(1'b1), .QN(n7539)
         );
  DFFSRX1 g4294_reg ( .D(n6580), .CK(clk), .RN(n8037), .SN(1'b1), .Q(g10122), 
        .QN(n5677) );
  DFFSRX1 g4300_reg ( .D(n6579), .CK(clk), .RN(n8058), .SN(1'b1), .Q(n12462)
         );
  DFFSRX1 g4311_reg ( .D(n6578), .CK(clk), .RN(n8028), .SN(1'b1), .Q(n7375), 
        .QN(n12541) );
  DFFSRX1 g4322_reg ( .D(n6577), .CK(clk), .RN(n8027), .SN(1'b1), .Q(n7252), 
        .QN(n12540) );
  DFFSRX1 g4332_reg ( .D(n6576), .CK(clk), .RN(n8027), .SN(1'b1), .Q(n7364), 
        .QN(n12539) );
  DFFSRX1 g4340_reg ( .D(n6575), .CK(clk), .RN(n8028), .SN(1'b1), .Q(n7412), 
        .QN(n12453) );
  DFFSRX1 g4349_reg ( .D(n6574), .CK(clk), .RN(n8028), .SN(1'b1), .Q(n7409), 
        .QN(n12452) );
  DFFSRX1 g4358_reg ( .D(n6573), .CK(clk), .RN(n8028), .SN(1'b1), .Q(n7353), 
        .QN(n12451) );
  DFFSRX1 g3990_reg ( .D(n6572), .CK(clk), .RN(n8031), .SN(1'b1), .Q(n12521), 
        .QN(n7542) );
  DFFSRX1 g4000_reg ( .D(n6571), .CK(clk), .RN(n8031), .SN(1'b1), .Q(g14518)
         );
  DFFSRX1 g4005_reg ( .D(n6570), .CK(clk), .RN(n8031), .SN(1'b1), .Q(g11418)
         );
  DFFSRX1 g4012_reg ( .D(n6569), .CK(clk), .RN(n8031), .SN(1'b1), .Q(g16775), 
        .QN(n5719) );
  DFFSRX1 g3969_reg ( .D(n6568), .CK(clk), .RN(n8031), .SN(1'b1), .Q(g16659), 
        .QN(n5720) );
  DFFSRX1 g3976_reg ( .D(g16659), .CK(clk), .RN(n8031), .SN(1'b1), .Q(g16693), 
        .QN(n7829) );
  DFFSRX1 g3983_reg ( .D(n6567), .CK(clk), .RN(n8031), .SN(1'b1), .Q(g13966)
         );
  DFFSRX1 g4027_reg ( .D(g13906), .CK(clk), .RN(n8031), .SN(1'b1), .Q(g16748)
         );
  DFFSRX1 g4031_reg ( .D(g16748), .CK(clk), .RN(n8030), .SN(1'b1), .Q(n12517)
         );
  DFFSRX1 g3639_reg ( .D(n6565), .CK(clk), .RN(n8064), .SN(1'b1), .Q(n12570), 
        .QN(n7543) );
  DFFSRX1 g3649_reg ( .D(n6564), .CK(clk), .RN(n8064), .SN(1'b1), .Q(g14451)
         );
  DFFSRX1 g3654_reg ( .D(n6563), .CK(clk), .RN(n8065), .SN(1'b1), .Q(g11388)
         );
  DFFSRX1 g3661_reg ( .D(n6562), .CK(clk), .RN(n8065), .SN(1'b1), .Q(g16744), 
        .QN(n5745) );
  DFFSRX1 g3618_reg ( .D(n6561), .CK(clk), .RN(n8065), .SN(1'b1), .Q(g16627), 
        .QN(n5746) );
  DFFSRX1 g3625_reg ( .D(g16627), .CK(clk), .RN(n8065), .SN(1'b1), .Q(g16656), 
        .QN(n7833) );
  DFFSRX1 g3632_reg ( .D(n6560), .CK(clk), .RN(n8065), .SN(1'b1), .Q(g13926)
         );
  DFFSRX1 g3676_reg ( .D(g13881), .CK(clk), .RN(n8064), .SN(1'b1), .Q(g16722)
         );
  DFFSRX1 g3680_reg ( .D(g16722), .CK(clk), .RN(n8064), .SN(1'b1), .Q(n12566)
         );
  DFFSRX1 g6682_reg ( .D(n6558), .CK(clk), .RN(n8037), .SN(1'b1), .Q(n12305), 
        .QN(n7544) );
  DFFSRX1 g6692_reg ( .D(n6557), .CK(clk), .RN(n8033), .SN(1'b1), .Q(g13099)
         );
  DFFSRX1 g6697_reg ( .D(n6556), .CK(clk), .RN(n8033), .SN(1'b1), .Q(g12470)
         );
  DFFSRX1 g6500_reg ( .D(n6555), .CK(clk), .RN(n8036), .SN(1'b1), .QN(n12183)
         );
  DFFSRX1 g6505_reg ( .D(n6554), .CK(clk), .RN(n8035), .SN(1'b1), .Q(n12184), 
        .QN(n7678) );
  DFFSRX1 g6509_reg ( .D(n6553), .CK(clk), .RN(n8036), .SN(1'b1), .Q(n12670), 
        .QN(n7318) );
  DFFSRX1 g6513_reg ( .D(n6552), .CK(clk), .RN(n8036), .SN(1'b1), .Q(n12176), 
        .QN(n7567) );
  DFFSRX1 g6519_reg ( .D(n6551), .CK(clk), .RN(n8032), .SN(1'b1), .QN(n7656)
         );
  DFFSRX1 g6523_reg ( .D(n6550), .CK(clk), .RN(n8036), .SN(1'b1), .Q(n12692), 
        .QN(n7579) );
  DFFSRX1 g6527_reg ( .D(n6549), .CK(clk), .RN(n8036), .SN(1'b1), .Q(n12175), 
        .QN(n7582) );
  DFFSRX1 g6533_reg ( .D(n6548), .CK(clk), .RN(n8035), .SN(1'b1), .Q(n12174)
         );
  DFFSRX1 g6537_reg ( .D(n6547), .CK(clk), .RN(n8036), .SN(1'b1), .Q(n12693), 
        .QN(n7323) );
  DFFSRX1 g6549_reg ( .D(n6546), .CK(clk), .RN(n8036), .SN(1'b1), .QN(n12173)
         );
  DFFSRX1 g6555_reg ( .D(n6545), .CK(clk), .RN(n8036), .SN(1'b1), .Q(n7426), 
        .QN(n12172) );
  DFFSRX1 g6561_reg ( .D(n6544), .CK(clk), .RN(n8036), .SN(1'b1), .Q(n12181), 
        .QN(n7260) );
  DFFSRX1 g6565_reg ( .D(n6543), .CK(clk), .RN(n8036), .SN(1'b1), .QN(n12182)
         );
  DFFSRX1 g6573_reg ( .D(n6542), .CK(clk), .RN(n8036), .SN(1'b1), .Q(n12185), 
        .QN(n7482) );
  DFFSRX1 g6581_reg ( .D(n6541), .CK(clk), .RN(n8035), .SN(1'b1), .Q(n12279)
         );
  DFFSRX1 g6605_reg ( .D(n6540), .CK(clk), .RN(n8035), .SN(1'b1), .Q(n12295)
         );
  DFFSRX1 g6609_reg ( .D(n6539), .CK(clk), .RN(n8035), .SN(1'b1), .Q(n12282)
         );
  DFFSRX1 g6625_reg ( .D(n6538), .CK(clk), .RN(n8035), .SN(1'b1), .Q(n12283)
         );
  DFFSRX1 g6641_reg ( .D(n6537), .CK(clk), .RN(n8035), .SN(1'b1), .Q(n12284)
         );
  DFFSRX1 g6589_reg ( .D(n6536), .CK(clk), .RN(n8035), .SN(1'b1), .Q(n12280)
         );
  DFFSRX1 g6585_reg ( .D(n6535), .CK(clk), .RN(n8035), .SN(1'b1), .Q(n7441), 
        .QN(n12281) );
  DFFSRX1 g6613_reg ( .D(n6534), .CK(clk), .RN(n8034), .SN(1'b1), .Q(n12291)
         );
  DFFSRX1 g6629_reg ( .D(n6533), .CK(clk), .RN(n8034), .SN(1'b1), .Q(n12292)
         );
  DFFSRX1 g6645_reg ( .D(n6532), .CK(clk), .RN(n8034), .SN(1'b1), .Q(n12290)
         );
  DFFSRX1 g6597_reg ( .D(n6531), .CK(clk), .RN(n8034), .SN(1'b1), .Q(n12285)
         );
  DFFSRX1 g6593_reg ( .D(n6530), .CK(clk), .RN(n8034), .SN(1'b1), .Q(n12293)
         );
  DFFSRX1 g6617_reg ( .D(n6529), .CK(clk), .RN(n8034), .SN(1'b1), .Q(n12296)
         );
  DFFSRX1 g6633_reg ( .D(n6528), .CK(clk), .RN(n8034), .SN(1'b1), .Q(n12297)
         );
  DFFSRX1 g6601_reg ( .D(n6527), .CK(clk), .RN(n8035), .SN(1'b1), .Q(n7388) );
  DFFSRX1 g6621_reg ( .D(n6526), .CK(clk), .RN(n8035), .SN(1'b1), .Q(n12289)
         );
  DFFSRX1 g6637_reg ( .D(n6525), .CK(clk), .RN(n8035), .SN(1'b1), .Q(n12287)
         );
  DFFSRX1 g6649_reg ( .D(n6524), .CK(clk), .RN(n8034), .SN(1'b1), .Q(n12286)
         );
  DFFSRX1 g6653_reg ( .D(n6523), .CK(clk), .RN(n8034), .SN(1'b1), .Q(n12288), 
        .QN(n7796) );
  DFFSRX1 g6657_reg ( .D(n6522), .CK(clk), .RN(n8034), .SN(1'b1), .Q(n12299)
         );
  DFFSRX1 g5016_reg ( .D(n6521), .CK(clk), .RN(n8029), .SN(1'b1), .Q(n7376), 
        .QN(n12276) );
  DFFSRX1 g5029_reg ( .D(n6520), .CK(clk), .RN(n8029), .SN(1'b1), .Q(n7270), 
        .QN(n12271) );
  DFFSRX1 g5033_reg ( .D(n6519), .CK(clk), .RN(n8029), .SN(1'b1), .Q(n12270), 
        .QN(n7399) );
  DFFSRX1 g5037_reg ( .D(n6518), .CK(clk), .RN(n8029), .SN(1'b1), .Q(n7427), 
        .QN(n12269) );
  DFFSRX1 g5041_reg ( .D(n6517), .CK(clk), .RN(n8029), .SN(1'b1), .Q(n12268), 
        .QN(n7408) );
  DFFSRX1 g5046_reg ( .D(n6516), .CK(clk), .RN(n8029), .SN(1'b1), .Q(n7358), 
        .QN(n12274) );
  DFFSRX1 g5052_reg ( .D(n6515), .CK(clk), .RN(n8029), .SN(1'b1), .QN(n12273)
         );
  DFFSRX1 g5057_reg ( .D(n6514), .CK(clk), .RN(n8028), .SN(1'b1), .QN(n12275)
         );
  DFFSRX1 g5062_reg ( .D(n6513), .CK(clk), .RN(n8030), .SN(1'b1), .Q(n12277), 
        .QN(n7406) );
  DFFSRX1 g5069_reg ( .D(n6512), .CK(clk), .RN(n8028), .SN(1'b1), .Q(n12265), 
        .QN(n7349) );
  DFFSRX1 g5073_reg ( .D(n6511), .CK(clk), .RN(n8030), .SN(1'b1), .Q(n12264), 
        .QN(n7750) );
  DFFSRX1 g5077_reg ( .D(n6510), .CK(clk), .RN(n8028), .SN(1'b1), .Q(n7327), 
        .QN(n12263) );
  DFFSRX1 g5084_reg ( .D(n6509), .CK(clk), .RN(n8030), .SN(1'b1), .Q(n7243) );
  DFFSRX1 g5080_reg ( .D(n6508), .CK(clk), .RN(n8030), .SN(1'b1), .QN(n12262)
         );
  DFFSRX1 g5092_reg ( .D(n6507), .CK(clk), .RN(n8030), .SN(1'b1), .Q(n12261), 
        .QN(n7471) );
  DFFSRX1 g5097_reg ( .D(n6506), .CK(clk), .RN(n8029), .SN(1'b1), .Q(n7498), 
        .QN(n12260) );
  DFFSRX1 g5101_reg ( .D(n6505), .CK(clk), .RN(n8029), .SN(1'b1), .Q(g9497), 
        .QN(n3814) );
  DFFSRX1 g5105_reg ( .D(n6504), .CK(clk), .RN(n8030), .SN(1'b1), .Q(g9553), 
        .QN(n3816) );
  DFFSRX1 g5115_reg ( .D(n6503), .CK(clk), .RN(n8028), .SN(1'b1), .QN(n12257)
         );
  DFFSRX1 g5124_reg ( .D(n6502), .CK(clk), .RN(n8074), .SN(1'b1), .QN(n7823)
         );
  DFFSRX1 g5128_reg ( .D(n6501), .CK(clk), .RN(n8074), .SN(1'b1), .Q(n12253), 
        .QN(n7568) );
  DFFSRX1 g5134_reg ( .D(n6500), .CK(clk), .RN(n8074), .SN(1'b1), .QN(n12252)
         );
  DFFSRX1 g5138_reg ( .D(n6499), .CK(clk), .RN(n8074), .SN(1'b1), .QN(n12694)
         );
  DFFSRX1 g5142_reg ( .D(n6498), .CK(clk), .RN(n8074), .SN(1'b1), .Q(n12251), 
        .QN(n7583) );
  DFFSRX1 g5148_reg ( .D(n6497), .CK(clk), .RN(n8073), .SN(1'b1), .Q(n12250)
         );
  DFFSRX1 g5152_reg ( .D(n6496), .CK(clk), .RN(n8074), .SN(1'b1), .QN(n7646)
         );
  DFFSRX1 g5164_reg ( .D(n6495), .CK(clk), .RN(n8074), .SN(1'b1), .QN(n12249)
         );
  DFFSRX1 g5170_reg ( .D(n6494), .CK(clk), .RN(n8073), .SN(1'b1), .Q(n7428), 
        .QN(n12248) );
  DFFSRX1 g5176_reg ( .D(n6493), .CK(clk), .RN(n8073), .SN(1'b1), .Q(n12255), 
        .QN(n7264) );
  DFFSRX1 g5180_reg ( .D(n6492), .CK(clk), .RN(n8073), .SN(1'b1), .QN(n12256)
         );
  DFFSRX1 g5188_reg ( .D(n6491), .CK(clk), .RN(n8073), .SN(1'b1), .Q(n12259), 
        .QN(n7493) );
  DFFSRX1 g5196_reg ( .D(n6490), .CK(clk), .RN(n8056), .SN(1'b1), .Q(n12975)
         );
  DFFSRX1 g5220_reg ( .D(n6489), .CK(clk), .RN(n8073), .SN(1'b1), .Q(n12981)
         );
  DFFSRX1 g5224_reg ( .D(n6488), .CK(clk), .RN(n8056), .SN(1'b1), .Q(n12977)
         );
  DFFSRX1 g5240_reg ( .D(n6487), .CK(clk), .RN(n8056), .SN(1'b1), .Q(n12978)
         );
  DFFSRX1 g5256_reg ( .D(n6486), .CK(clk), .RN(n8056), .SN(1'b1), .Q(n7227) );
  DFFSRX1 g5204_reg ( .D(n6485), .CK(clk), .RN(n8052), .SN(1'b1), .Q(n12976)
         );
  DFFSRX1 g5200_reg ( .D(n6484), .CK(clk), .RN(n8052), .SN(1'b1), .Q(n7446), 
        .QN(n12974) );
  DFFSRX1 g5228_reg ( .D(n6483), .CK(clk), .RN(n8052), .SN(1'b1), .Q(n12987)
         );
  DFFSRX1 g5244_reg ( .D(n6482), .CK(clk), .RN(n8052), .SN(1'b1), .Q(n12986)
         );
  DFFSRX1 g5260_reg ( .D(n6481), .CK(clk), .RN(n8052), .SN(1'b1), .Q(n12988)
         );
  DFFSRX1 g5212_reg ( .D(n6480), .CK(clk), .RN(n8051), .SN(1'b1), .Q(n12989)
         );
  DFFSRX1 g5208_reg ( .D(n6479), .CK(clk), .RN(n8051), .SN(1'b1), .Q(n12979)
         );
  DFFSRX1 g5232_reg ( .D(n6478), .CK(clk), .RN(n8051), .SN(1'b1), .Q(n12994)
         );
  DFFSRX1 g5248_reg ( .D(n6477), .CK(clk), .RN(n8051), .SN(1'b1), .Q(n12991)
         );
  DFFSRX1 g5216_reg ( .D(n6476), .CK(clk), .RN(n8073), .SN(1'b1), .Q(n12985)
         );
  DFFSRX1 g5236_reg ( .D(n6475), .CK(clk), .RN(n8073), .SN(1'b1), .Q(n12982)
         );
  DFFSRX1 g5252_reg ( .D(n6474), .CK(clk), .RN(n8073), .SN(1'b1), .Q(n12983)
         );
  DFFSRX1 g5264_reg ( .D(n6473), .CK(clk), .RN(n8051), .SN(1'b1), .Q(n12990)
         );
  DFFSRX1 g5268_reg ( .D(n6472), .CK(clk), .RN(n8073), .SN(1'b1), .Q(n12984), 
        .QN(n7798) );
  DFFSRX1 g5272_reg ( .D(n6471), .CK(clk), .RN(n8073), .SN(1'b1), .Q(n13005)
         );
  DFFSRX1 g5276_reg ( .D(n6470), .CK(clk), .RN(n8073), .SN(1'b1), .Q(g17519), 
        .QN(n5604) );
  DFFSRX1 g5283_reg ( .D(g17519), .CK(clk), .RN(n8072), .SN(1'b1), .Q(g17577), 
        .QN(n7821) );
  DFFSRX1 g5313_reg ( .D(n6469), .CK(clk), .RN(n8072), .SN(1'b1), .Q(g12238)
         );
  DFFSRX1 g5290_reg ( .D(n6468), .CK(clk), .RN(n8072), .SN(1'b1), .Q(g14662)
         );
  DFFSRX1 g5320_reg ( .D(n6467), .CK(clk), .RN(n8072), .SN(1'b1), .Q(g17674), 
        .QN(n5605) );
  DFFSRX1 g5335_reg ( .D(g14597), .CK(clk), .RN(n8071), .SN(1'b1), .Q(g17639)
         );
  DFFSRX1 g5339_reg ( .D(g17639), .CK(clk), .RN(n8071), .SN(1'b1), .Q(n12980), 
        .QN(n7799) );
  DFFSRX1 g5343_reg ( .D(n6465), .CK(clk), .RN(n8072), .SN(1'b1), .Q(g25219), 
        .QN(n302) );
  DFFSRX1 g5348_reg ( .D(n6464), .CK(clk), .RN(n8072), .SN(1'b1), .QN(n7657)
         );
  DFFSRX1 g5352_reg ( .D(n6463), .CK(clk), .RN(n8072), .SN(1'b1), .Q(n12384), 
        .QN(n7626) );
  DFFSRX1 g5357_reg ( .D(n6462), .CK(clk), .RN(n8072), .SN(1'b1), .Q(n7366), 
        .QN(n12992) );
  DFFSRX1 g5448_reg ( .D(n6461), .CK(clk), .RN(n8040), .SN(1'b1), .Q(g9555), 
        .QN(n7990) );
  DFFSRX1 g5452_reg ( .D(n6460), .CK(clk), .RN(n8040), .SN(1'b1), .Q(g9615), 
        .QN(n3818) );
  DFFSRX1 g5297_reg ( .D(n6459), .CK(clk), .RN(n8072), .SN(1'b1), .Q(n12993)
         );
  DFFSRX1 g4704_reg ( .D(n6458), .CK(clk), .RN(n8071), .SN(1'b1), .Q(n7459) );
  DFFSRX1 g4709_reg ( .D(n6457), .CK(clk), .RN(n8071), .SN(1'b1), .Q(n7380), 
        .QN(n13004) );
  DFFSRX1 g4717_reg ( .D(n6456), .CK(clk), .RN(n8071), .SN(1'b1), .Q(n12398)
         );
  DFFSRX1 g4722_reg ( .D(n6455), .CK(clk), .RN(n8071), .SN(1'b1), .Q(n12397)
         );
  DFFSRX1 g4737_reg ( .D(n6454), .CK(clk), .RN(n8071), .SN(1'b1), .Q(n12399), 
        .QN(n7751) );
  DFFSRX1 g4743_reg ( .D(n6453), .CK(clk), .RN(n8071), .SN(1'b1), .Q(n7442), 
        .QN(n12401) );
  DFFSRX1 g4749_reg ( .D(n6452), .CK(clk), .RN(n8071), .SN(1'b1), .Q(n12383), 
        .QN(n7780) );
  DFFSRX1 g4776_reg ( .D(n6451), .CK(clk), .RN(n8045), .SN(1'b1), .Q(n7246), 
        .QN(n13001) );
  DFFSRX1 g4785_reg ( .D(n6450), .CK(clk), .RN(n8045), .SN(1'b1), .Q(n7249), 
        .QN(n13003) );
  DFFSRX1 g4793_reg ( .D(n6449), .CK(clk), .RN(n8045), .SN(1'b1), .Q(n7354), 
        .QN(n13000) );
  DFFSRX1 g4801_reg ( .D(n6448), .CK(clk), .RN(n8045), .SN(1'b1), .Q(n7255), 
        .QN(n12997) );
  DFFSRX1 g5808_reg ( .D(n6447), .CK(clk), .RN(n8030), .SN(1'b1), .QN(n12212)
         );
  DFFSRX1 g5821_reg ( .D(n6446), .CK(clk), .RN(n8071), .SN(1'b1), .Q(n12208), 
        .QN(n7569) );
  DFFSRX1 g5827_reg ( .D(n6445), .CK(clk), .RN(n8053), .SN(1'b1), .QN(n12207)
         );
  DFFSRX1 g5831_reg ( .D(n6444), .CK(clk), .RN(n8070), .SN(1'b1), .QN(n12691)
         );
  DFFSRX1 g5835_reg ( .D(n6443), .CK(clk), .RN(n8070), .SN(1'b1), .Q(n12206), 
        .QN(n7584) );
  DFFSRX1 g5841_reg ( .D(n6442), .CK(clk), .RN(n8070), .SN(1'b1), .Q(n12205)
         );
  DFFSRX1 g5845_reg ( .D(n6441), .CK(clk), .RN(n8070), .SN(1'b1), .QN(n7641)
         );
  DFFSRX1 g5857_reg ( .D(n6440), .CK(clk), .RN(n8070), .SN(1'b1), .QN(n12204)
         );
  DFFSRX1 g5863_reg ( .D(n6439), .CK(clk), .RN(n8070), .SN(1'b1), .Q(n7429), 
        .QN(n12203) );
  DFFSRX1 g5869_reg ( .D(n6438), .CK(clk), .RN(n8070), .SN(1'b1), .Q(n12210), 
        .QN(n7261) );
  DFFSRX1 g5873_reg ( .D(n6437), .CK(clk), .RN(n8070), .SN(1'b1), .QN(n12211)
         );
  DFFSRX1 g5881_reg ( .D(n6436), .CK(clk), .RN(n8070), .SN(1'b1), .Q(n12214), 
        .QN(n7483) );
  DFFSRX1 g5889_reg ( .D(n6435), .CK(clk), .RN(n8056), .SN(1'b1), .Q(n12313)
         );
  DFFSRX1 g5913_reg ( .D(n6434), .CK(clk), .RN(n8070), .SN(1'b1), .Q(n12310)
         );
  DFFSRX1 g5917_reg ( .D(n6433), .CK(clk), .RN(n8056), .SN(1'b1), .Q(n12323)
         );
  DFFSRX1 g5933_reg ( .D(n6432), .CK(clk), .RN(n8054), .SN(1'b1), .Q(n12324)
         );
  DFFSRX1 g5949_reg ( .D(n6431), .CK(clk), .RN(n8054), .SN(1'b1), .Q(n12325)
         );
  DFFSRX1 g5897_reg ( .D(n6430), .CK(clk), .RN(n8054), .SN(1'b1), .Q(n12314)
         );
  DFFSRX1 g5893_reg ( .D(n6429), .CK(clk), .RN(n8055), .SN(1'b1), .Q(n7443), 
        .QN(n12316) );
  DFFSRX1 g5921_reg ( .D(n6428), .CK(clk), .RN(n8054), .SN(1'b1), .Q(n12318)
         );
  DFFSRX1 g5937_reg ( .D(n6427), .CK(clk), .RN(n8054), .SN(1'b1), .Q(n12319)
         );
  DFFSRX1 g5953_reg ( .D(n6426), .CK(clk), .RN(n8054), .SN(1'b1), .Q(n12317)
         );
  DFFSRX1 g5905_reg ( .D(n6425), .CK(clk), .RN(n8054), .SN(1'b1), .Q(n12307)
         );
  DFFSRX1 g5901_reg ( .D(n6424), .CK(clk), .RN(n8054), .SN(1'b1), .Q(n12309)
         );
  DFFSRX1 g5925_reg ( .D(n6423), .CK(clk), .RN(n8054), .SN(1'b1), .Q(n12311)
         );
  DFFSRX1 g5941_reg ( .D(n6422), .CK(clk), .RN(n8054), .SN(1'b1), .Q(n12312)
         );
  DFFSRX1 g5909_reg ( .D(n6421), .CK(clk), .RN(n8070), .SN(1'b1), .Q(n7389) );
  DFFSRX1 g5929_reg ( .D(n6420), .CK(clk), .RN(n8054), .SN(1'b1), .Q(n12322)
         );
  DFFSRX1 g5945_reg ( .D(n6419), .CK(clk), .RN(n8054), .SN(1'b1), .Q(n12320)
         );
  DFFSRX1 g5957_reg ( .D(n6418), .CK(clk), .RN(n8053), .SN(1'b1), .Q(n12308)
         );
  DFFSRX1 g5961_reg ( .D(n6417), .CK(clk), .RN(n8053), .SN(1'b1), .Q(n12321), 
        .QN(n7802) );
  DFFSRX1 g5965_reg ( .D(n6416), .CK(clk), .RN(n8053), .SN(1'b1), .Q(n12327)
         );
  DFFSRX1 g5969_reg ( .D(n6415), .CK(clk), .RN(n8053), .SN(1'b1), .Q(g17607), 
        .QN(n5568) );
  DFFSRX1 g5976_reg ( .D(g17607), .CK(clk), .RN(n8053), .SN(1'b1), .Q(g17646), 
        .QN(n7813) );
  DFFSRX1 g6005_reg ( .D(n6414), .CK(clk), .RN(n8052), .SN(1'b1), .Q(g12350)
         );
  DFFSRX1 g5983_reg ( .D(n6413), .CK(clk), .RN(n8052), .SN(1'b1), .Q(g14738)
         );
  DFFSRX1 g6012_reg ( .D(n6412), .CK(clk), .RN(n8052), .SN(1'b1), .Q(g17739), 
        .QN(n5569) );
  DFFSRX1 g6027_reg ( .D(g14673), .CK(clk), .RN(n8052), .SN(1'b1), .Q(g17715), 
        .QN(n7618) );
  DFFSRX1 g6031_reg ( .D(g17715), .CK(clk), .RN(n8052), .SN(1'b1), .Q(n12315), 
        .QN(n7803) );
  DFFSRX1 g6035_reg ( .D(n6411), .CK(clk), .RN(n8053), .SN(1'b1), .Q(n7416), 
        .QN(n12326) );
  DFFSRX1 g5798_reg ( .D(n6410), .CK(clk), .RN(n8040), .SN(1'b1), .Q(g9680), 
        .QN(n3820) );
  DFFSRX1 g5794_reg ( .D(n6409), .CK(clk), .RN(n8040), .SN(1'b1), .Q(g9617), 
        .QN(n7992) );
  DFFSRX1 g6040_reg ( .D(n6408), .CK(clk), .RN(n8053), .SN(1'b1), .QN(n7659)
         );
  DFFSRX1 g6044_reg ( .D(n6407), .CK(clk), .RN(n8053), .SN(1'b1), .Q(n12376)
         );
  DFFSRX1 g6049_reg ( .D(n6406), .CK(clk), .RN(n8053), .SN(1'b1), .Q(n7253), 
        .QN(n12378) );
  DFFSRX1 g5990_reg ( .D(n6405), .CK(clk), .RN(n8053), .SN(1'b1), .Q(n12377), 
        .QN(n7547) );
  DFFSRX1 g6000_reg ( .D(n6404), .CK(clk), .RN(n8053), .SN(1'b1), .Q(g13068)
         );
  DFFSRX1 g6154_reg ( .D(n6403), .CK(clk), .RN(n8038), .SN(1'b1), .QN(n12198)
         );
  DFFSRX1 g6167_reg ( .D(n6402), .CK(clk), .RN(n8038), .SN(1'b1), .Q(n12194), 
        .QN(n7570) );
  DFFSRX1 g6173_reg ( .D(n6401), .CK(clk), .RN(n8038), .SN(1'b1), .QN(n12193)
         );
  DFFSRX1 g6177_reg ( .D(n6400), .CK(clk), .RN(n8038), .SN(1'b1), .QN(n12690)
         );
  DFFSRX1 g6181_reg ( .D(n6399), .CK(clk), .RN(n8038), .SN(1'b1), .Q(n12192), 
        .QN(n7585) );
  DFFSRX1 g6187_reg ( .D(n6398), .CK(clk), .RN(n8038), .SN(1'b1), .Q(n12191)
         );
  DFFSRX1 g6191_reg ( .D(n6397), .CK(clk), .RN(n8037), .SN(1'b1), .QN(n7642)
         );
  DFFSRX1 g6203_reg ( .D(n6396), .CK(clk), .RN(n8047), .SN(1'b1), .QN(n12190)
         );
  DFFSRX1 g6209_reg ( .D(n6395), .CK(clk), .RN(n8047), .SN(1'b1), .Q(n7430), 
        .QN(n12189) );
  DFFSRX1 g6215_reg ( .D(n6394), .CK(clk), .RN(n8047), .SN(1'b1), .Q(n12196), 
        .QN(n7262) );
  DFFSRX1 g6219_reg ( .D(n6393), .CK(clk), .RN(n8047), .SN(1'b1), .QN(n12197)
         );
  DFFSRX1 g6227_reg ( .D(n6392), .CK(clk), .RN(n8047), .SN(1'b1), .Q(n12200), 
        .QN(n7484) );
  DFFSRX1 g6235_reg ( .D(n6391), .CK(clk), .RN(n8047), .SN(1'b1), .Q(n12336)
         );
  DFFSRX1 g6259_reg ( .D(n6390), .CK(clk), .RN(n8047), .SN(1'b1), .Q(n12333)
         );
  DFFSRX1 g6263_reg ( .D(n6389), .CK(clk), .RN(n8047), .SN(1'b1), .Q(n12346)
         );
  DFFSRX1 g6279_reg ( .D(n6388), .CK(clk), .RN(n8047), .SN(1'b1), .Q(n12347)
         );
  DFFSRX1 g6295_reg ( .D(n6387), .CK(clk), .RN(n8046), .SN(1'b1), .Q(n12348)
         );
  DFFSRX1 g6243_reg ( .D(n6386), .CK(clk), .RN(n8046), .SN(1'b1), .Q(n12337)
         );
  DFFSRX1 g6239_reg ( .D(n6385), .CK(clk), .RN(n8046), .SN(1'b1), .Q(n7444), 
        .QN(n12339) );
  DFFSRX1 g6267_reg ( .D(n6384), .CK(clk), .RN(n8046), .SN(1'b1), .Q(n12341)
         );
  DFFSRX1 g6283_reg ( .D(n6383), .CK(clk), .RN(n8046), .SN(1'b1), .Q(n12342)
         );
  DFFSRX1 g6299_reg ( .D(n6382), .CK(clk), .RN(n8046), .SN(1'b1), .Q(n12340)
         );
  DFFSRX1 g6251_reg ( .D(n6381), .CK(clk), .RN(n8046), .SN(1'b1), .Q(n12330)
         );
  DFFSRX1 g6247_reg ( .D(n6380), .CK(clk), .RN(n8046), .SN(1'b1), .Q(n12332)
         );
  DFFSRX1 g6271_reg ( .D(n6379), .CK(clk), .RN(n8046), .SN(1'b1), .Q(n12334)
         );
  DFFSRX1 g6287_reg ( .D(n6378), .CK(clk), .RN(n8046), .SN(1'b1), .Q(n12335)
         );
  DFFSRX1 g6255_reg ( .D(n6377), .CK(clk), .RN(n8047), .SN(1'b1), .Q(n7390) );
  DFFSRX1 g6275_reg ( .D(n6376), .CK(clk), .RN(n8047), .SN(1'b1), .Q(n12345)
         );
  DFFSRX1 g6291_reg ( .D(n6375), .CK(clk), .RN(n8047), .SN(1'b1), .Q(n12343)
         );
  DFFSRX1 g6303_reg ( .D(n6374), .CK(clk), .RN(n8046), .SN(1'b1), .Q(n12331)
         );
  DFFSRX1 g6307_reg ( .D(n6373), .CK(clk), .RN(n8046), .SN(1'b1), .Q(n12344), 
        .QN(n7804) );
  DFFSRX1 g6311_reg ( .D(n6372), .CK(clk), .RN(n8045), .SN(1'b1), .Q(n12350)
         );
  DFFSRX1 g6315_reg ( .D(n6371), .CK(clk), .RN(n8045), .SN(1'b1), .Q(g17649), 
        .QN(n5537) );
  DFFSRX1 g6322_reg ( .D(g17649), .CK(clk), .RN(n8045), .SN(1'b1), .Q(g17685), 
        .QN(n7809) );
  DFFSRX1 g6351_reg ( .D(n6370), .CK(clk), .RN(n8044), .SN(1'b1), .Q(g12422)
         );
  DFFSRX1 g6329_reg ( .D(n6369), .CK(clk), .RN(n8044), .SN(1'b1), .Q(g14779)
         );
  DFFSRX1 g6358_reg ( .D(n6368), .CK(clk), .RN(n8044), .SN(1'b1), .Q(g17760), 
        .QN(n5538) );
  DFFSRX1 g6373_reg ( .D(g14705), .CK(clk), .RN(n8044), .SN(1'b1), .Q(g17743), 
        .QN(n7596) );
  DFFSRX1 g6377_reg ( .D(g17743), .CK(clk), .RN(n8044), .SN(1'b1), .Q(n12338), 
        .QN(n7806) );
  DFFSRX1 g6381_reg ( .D(n6367), .CK(clk), .RN(n8045), .SN(1'b1), .Q(n7417), 
        .QN(n12349) );
  DFFSRX1 g6144_reg ( .D(n6366), .CK(clk), .RN(n8039), .SN(1'b1), .Q(g9741), 
        .QN(n3822) );
  DFFSRX1 g6140_reg ( .D(n6365), .CK(clk), .RN(n8038), .SN(1'b1), .Q(g9682), 
        .QN(n7994) );
  DFFSRX1 g6386_reg ( .D(n6364), .CK(clk), .RN(n8045), .SN(1'b1), .QN(n7660)
         );
  DFFSRX1 g6390_reg ( .D(n6363), .CK(clk), .RN(n8045), .SN(1'b1), .Q(n12372)
         );
  DFFSRX1 g6395_reg ( .D(n6362), .CK(clk), .RN(n8044), .SN(1'b1), .Q(n7254), 
        .QN(n12374) );
  DFFSRX1 g6336_reg ( .D(n6361), .CK(clk), .RN(n8044), .SN(1'b1), .Q(n12373), 
        .QN(n7548) );
  DFFSRX1 g6346_reg ( .D(n6360), .CK(clk), .RN(n8044), .SN(1'b1), .Q(g13085)
         );
  DFFSRX1 g4698_reg ( .D(n6359), .CK(clk), .RN(n8045), .SN(1'b1), .Q(n13002), 
        .QN(n7714) );
  DFFSRX1 g5308_reg ( .D(n6358), .CK(clk), .RN(n8072), .SN(1'b1), .Q(g13039)
         );
  DFFSRX1 g86_reg ( .D(n6357), .CK(clk), .RN(n8025), .SN(1'b1), .Q(g20557), 
        .QN(n5532) );
  DFFSRX1 g1227_reg ( .D(n6356), .CK(clk), .RN(n8020), .SN(1'b1), .Q(g12919), 
        .QN(n5888) );
  DFFSRX1 g1242_reg ( .D(n6355), .CK(clk), .RN(n8018), .SN(1'b1), .Q(g30332), 
        .QN(n5529) );
  DFFSRX1 g1246_reg ( .D(n6354), .CK(clk), .RN(n8018), .SN(1'b1), .Q(n7500), 
        .QN(n13006) );
  DFFSRX1 g1233_reg ( .D(n6353), .CK(clk), .RN(n8021), .SN(1'b1), .Q(g10500)
         );
  DFFSRX1 g1236_reg ( .D(g10500), .CK(clk), .RN(n8021), .SN(1'b1), .Q(n13062)
         );
  DFFSRX1 g996_reg ( .D(n6352), .CK(clk), .RN(n8020), .SN(1'b1), .Q(n13070), 
        .QN(n7494) );
  DFFSRX1 g1157_reg ( .D(n6351), .CK(clk), .RN(n8021), .SN(1'b1), .Q(g7916), 
        .QN(n763) );
  DFFSRX1 g1239_reg ( .D(n6350), .CK(clk), .RN(n8021), .SN(1'b1), .Q(g8416), 
        .QN(n5530) );
  DFFSRX1 g990_reg ( .D(n6349), .CK(clk), .RN(n8021), .SN(1'b1), .Q(n13075), 
        .QN(n7517) );
  DFFSRX1 g1036_reg ( .D(n6348), .CK(clk), .RN(n8019), .SN(1'b1), .Q(n13065)
         );
  DFFSRX1 g1041_reg ( .D(n6347), .CK(clk), .RN(n8019), .SN(1'b1), .Q(n13064), 
        .QN(n7715) );
  DFFSRX1 g1046_reg ( .D(n6346), .CK(clk), .RN(n8019), .SN(1'b1), .Q(n7445), 
        .QN(n13069) );
  DFFSRX1 g1008_reg ( .D(n6345), .CK(clk), .RN(n8020), .SN(1'b1), .Q(n13071), 
        .QN(n7382) );
  DFFSRX1 g1018_reg ( .D(n6344), .CK(clk), .RN(n8019), .SN(1'b1), .Q(n7418), 
        .QN(n13072) );
  DFFSRX1 g1024_reg ( .D(n6343), .CK(clk), .RN(n8019), .SN(1'b1), .Q(n13067), 
        .QN(n7571) );
  DFFSRX1 g1030_reg ( .D(n6342), .CK(clk), .RN(n8020), .SN(1'b1), .Q(n13073), 
        .QN(n7472) );
  DFFSRX1 g1002_reg ( .D(n6341), .CK(clk), .RN(n8020), .SN(1'b1), .Q(n13076), 
        .QN(n7476) );
  DFFSRX1 g1052_reg ( .D(n6340), .CK(clk), .RN(n8019), .SN(1'b1), .Q(n13063), 
        .QN(n7610) );
  DFFSRX1 g1056_reg ( .D(n6339), .CK(clk), .RN(n8019), .SN(1'b1), .Q(g19334), 
        .QN(n766) );
  DFFSRX1 g1061_reg ( .D(n6338), .CK(clk), .RN(n8022), .SN(1'b1), .Q(n13061), 
        .QN(n7533) );
  DFFSRX1 g1189_reg ( .D(n6337), .CK(clk), .RN(n8021), .SN(1'b1), .Q(n13055), 
        .QN(n7752) );
  DFFSRX1 g1193_reg ( .D(n6336), .CK(clk), .RN(n8020), .SN(1'b1), .Q(n13050), 
        .QN(n7690) );
  DFFSRX1 g1171_reg ( .D(n6335), .CK(clk), .RN(n8019), .SN(1'b1), .Q(n13053)
         );
  DFFSRX1 g1183_reg ( .D(n6334), .CK(clk), .RN(n8019), .SN(1'b1), .Q(n13054), 
        .QN(n7557) );
  DFFSRX1 g1178_reg ( .D(n6333), .CK(clk), .RN(n8019), .SN(1'b1), .Q(n13056), 
        .QN(n7635) );
  DFFSRX1 g1199_reg ( .D(n6332), .CK(clk), .RN(n8020), .SN(1'b1), .Q(n13052), 
        .QN(n7518) );
  DFFSRX1 g1070_reg ( .D(n6331), .CK(clk), .RN(n8021), .SN(1'b1), .Q(n13051), 
        .QN(n7628) );
  DFFSRX1 g1205_reg ( .D(n6330), .CK(clk), .RN(n8020), .SN(1'b1), .Q(n13047), 
        .QN(n7532) );
  DFFSRX1 g1211_reg ( .D(n6329), .CK(clk), .RN(n8020), .SN(1'b1), .Q(n13049), 
        .QN(n7537) );
  DFFSRX1 g1216_reg ( .D(n6328), .CK(clk), .RN(n8020), .SN(1'b1), .Q(n13016), 
        .QN(n7636) );
  DFFSRX1 g1221_reg ( .D(n6327), .CK(clk), .RN(n8020), .SN(1'b1), .Q(n13046), 
        .QN(n7549) );
  DFFSRX1 g1079_reg ( .D(g17291), .CK(clk), .RN(n8021), .SN(1'b1), .Q(g17316), 
        .QN(n7912) );
  DFFSRX1 g1083_reg ( .D(g17316), .CK(clk), .RN(n8021), .SN(1'b1), .Q(g17400), 
        .QN(n7933) );
  DFFSRX1 g1094_reg ( .D(n6326), .CK(clk), .RN(n8018), .SN(1'b1), .Q(n13044), 
        .QN(n7716) );
  DFFSRX1 g1099_reg ( .D(n6325), .CK(clk), .RN(n8018), .SN(1'b1), .Q(n13045), 
        .QN(n7272) );
  DFFSRX1 g1146_reg ( .D(n6324), .CK(clk), .RN(n8022), .SN(1'b1), .Q(n13043), 
        .QN(n7679) );
  DFFSRX1 g1152_reg ( .D(n6323), .CK(clk), .RN(n8019), .SN(1'b1), .Q(n13040), 
        .QN(n7371) );
  DFFSRX1 g1105_reg ( .D(n6322), .CK(clk), .RN(n8018), .SN(1'b1), .Q(n13038), 
        .QN(n7367) );
  DFFSRX1 g1124_reg ( .D(n6321), .CK(clk), .RN(n8018), .SN(1'b1), .Q(n13037), 
        .QN(n7807) );
  DFFSRX1 g1129_reg ( .D(n6320), .CK(clk), .RN(n8018), .SN(1'b1), .Q(n13036), 
        .QN(n7282) );
  DFFSRX1 g1135_reg ( .D(n6319), .CK(clk), .RN(n8018), .SN(1'b1), .Q(n13041), 
        .QN(n7356) );
  DFFSRX1 g1116_reg ( .D(n6318), .CK(clk), .RN(n8022), .SN(1'b1), .Q(g13259), 
        .QN(n768) );
  DFFSRX1 g1570_reg ( .D(n6317), .CK(clk), .RN(n8016), .SN(1'b1), .Q(g12923), 
        .QN(n5511) );
  DFFSRX1 g1585_reg ( .D(n6316), .CK(clk), .RN(n8014), .SN(1'b1), .Q(n12893), 
        .QN(n7474) );
  DFFSRX1 g1589_reg ( .D(n6315), .CK(clk), .RN(n8014), .SN(1'b1), .Q(n12895), 
        .QN(n7529) );
  DFFSRX1 g1576_reg ( .D(n6314), .CK(clk), .RN(n8017), .SN(1'b1), .Q(g10527)
         );
  DFFSRX1 g1579_reg ( .D(g10527), .CK(clk), .RN(n8017), .SN(1'b1), .Q(n12951)
         );
  DFFSRX1 g1582_reg ( .D(n6313), .CK(clk), .RN(n8017), .SN(1'b1), .Q(g8475) );
  DFFSRX1 g1333_reg ( .D(n6312), .CK(clk), .RN(n8017), .SN(1'b1), .Q(n12963), 
        .QN(n7478) );
  DFFSRX1 g1339_reg ( .D(n6311), .CK(clk), .RN(n8016), .SN(1'b1), .Q(n12966), 
        .QN(n7495) );
  DFFSRX1 g1500_reg ( .D(n6310), .CK(clk), .RN(n8017), .SN(1'b1), .Q(g7946), 
        .QN(n716) );
  DFFSRX1 g1532_reg ( .D(n6309), .CK(clk), .RN(n8015), .SN(1'b1), .Q(n12948), 
        .QN(n7753) );
  DFFSRX1 g1536_reg ( .D(n6308), .CK(clk), .RN(n8016), .SN(1'b1), .Q(n12945), 
        .QN(n7689) );
  DFFSRX1 g1542_reg ( .D(n6307), .CK(clk), .RN(n8016), .SN(1'b1), .Q(n12947), 
        .QN(n7519) );
  DFFSRX1 g1548_reg ( .D(n6306), .CK(clk), .RN(n8016), .SN(1'b1), .Q(n12942), 
        .QN(n7527) );
  DFFSRX1 g1554_reg ( .D(n6305), .CK(clk), .RN(n8016), .SN(1'b1), .Q(n12944), 
        .QN(n7509) );
  DFFSRX1 g1559_reg ( .D(n6304), .CK(clk), .RN(n8016), .SN(1'b1), .Q(n12897), 
        .QN(n7637) );
  DFFSRX1 g1564_reg ( .D(n6303), .CK(clk), .RN(n8016), .SN(1'b1), .Q(n7496), 
        .QN(n12941) );
  DFFSRX1 g1422_reg ( .D(g17320), .CK(clk), .RN(n8017), .SN(1'b1), .Q(g17404), 
        .QN(n7911) );
  DFFSRX1 g1426_reg ( .D(g17404), .CK(clk), .RN(n8017), .SN(1'b1), .Q(g17423), 
        .QN(n699) );
  DFFSRX1 g1430_reg ( .D(g17423), .CK(clk), .RN(n8017), .SN(1'b1), .Q(n12943), 
        .QN(n7313) );
  DFFSRX1 g1437_reg ( .D(n6302), .CK(clk), .RN(n8014), .SN(1'b1), .Q(n12912)
         );
  DFFSRX1 g1442_reg ( .D(n6301), .CK(clk), .RN(n8014), .SN(1'b1), .Q(n12971)
         );
  DFFSRX1 g1489_reg ( .D(n6300), .CK(clk), .RN(n8014), .SN(1'b1), .Q(n12911)
         );
  DFFSRX1 g1495_reg ( .D(n6299), .CK(clk), .RN(n8014), .SN(1'b1), .Q(n12969), 
        .QN(n7372) );
  DFFSRX1 g1300_reg ( .D(n6298), .CK(clk), .RN(n8018), .SN(1'b1), .Q(n12968), 
        .QN(n7534) );
  DFFSRX1 g1306_reg ( .D(n6297), .CK(clk), .RN(n8018), .SN(1'b1), .Q(n12965), 
        .QN(n7332) );
  DFFSRX1 g1312_reg ( .D(n6296), .CK(clk), .RN(n8018), .SN(1'b1), .Q(n12955), 
        .QN(n7612) );
  DFFSRX1 g1319_reg ( .D(n6295), .CK(clk), .RN(n8017), .SN(1'b1), .Q(n12952)
         );
  DFFSRX1 g1322_reg ( .D(n6294), .CK(clk), .RN(n8016), .SN(1'b1), .Q(n12964), 
        .QN(n7256) );
  DFFSRX1 g1379_reg ( .D(n6293), .CK(clk), .RN(n8015), .SN(1'b1), .Q(n12961)
         );
  DFFSRX1 g1384_reg ( .D(n6292), .CK(clk), .RN(n8015), .SN(1'b1), .Q(n12949), 
        .QN(n7718) );
  DFFSRX1 g1389_reg ( .D(n6291), .CK(clk), .RN(n8017), .SN(1'b1), .Q(n7501), 
        .QN(n12957) );
  DFFSRX1 g1351_reg ( .D(n6290), .CK(clk), .RN(n8015), .SN(1'b1), .Q(n12956), 
        .QN(n7383) );
  DFFSRX1 g1345_reg ( .D(n6289), .CK(clk), .RN(n8015), .SN(1'b1), .Q(n12962), 
        .QN(n7477) );
  DFFSRX1 g1361_reg ( .D(n6288), .CK(clk), .RN(n8015), .SN(1'b1), .Q(n7419), 
        .QN(n12958) );
  DFFSRX1 g1367_reg ( .D(n6287), .CK(clk), .RN(n8015), .SN(1'b1), .Q(n12960), 
        .QN(n7572) );
  DFFSRX1 g1373_reg ( .D(n6286), .CK(clk), .RN(n8015), .SN(1'b1), .Q(n12959), 
        .QN(n7473) );
  DFFSRX1 g1514_reg ( .D(n6285), .CK(clk), .RN(n8015), .SN(1'b1), .Q(n12973)
         );
  DFFSRX1 g1526_reg ( .D(n6284), .CK(clk), .RN(n8015), .SN(1'b1), .Q(n12972), 
        .QN(n7551) );
  DFFSRX1 g1521_reg ( .D(n6283), .CK(clk), .RN(n8015), .SN(1'b1), .Q(n12967), 
        .QN(n7638) );
  DFFSRX1 g1395_reg ( .D(n6282), .CK(clk), .RN(n8017), .SN(1'b1), .Q(n12953), 
        .QN(n7423) );
  DFFSRX1 g1399_reg ( .D(n6281), .CK(clk), .RN(n8015), .SN(1'b1), .Q(g19357), 
        .QN(n719) );
  DFFSRX1 g1459_reg ( .D(n6280), .CK(clk), .RN(n8016), .SN(1'b1), .Q(g13272), 
        .QN(n721) );
  DFFSRX1 g1467_reg ( .D(n6279), .CK(clk), .RN(n8014), .SN(1'b1), .Q(n12907), 
        .QN(n7808) );
  DFFSRX1 g1472_reg ( .D(n6278), .CK(clk), .RN(n8014), .SN(1'b1), .Q(n12908)
         );
  DFFSRX1 g1478_reg ( .D(n6277), .CK(clk), .RN(n8014), .SN(1'b1), .Q(n12913)
         );
  DFFSRX1 g1448_reg ( .D(n6276), .CK(clk), .RN(n8014), .SN(1'b1), .Q(n12909)
         );
  DFFSRX1 g1404_reg ( .D(n6275), .CK(clk), .RN(n8016), .SN(1'b1), .Q(n12954), 
        .QN(n7479) );
  DFFSRX1 g1413_reg ( .D(n6274), .CK(clk), .RN(n8016), .SN(1'b1), .Q(n12946), 
        .QN(n7629) );
  DFFSRX1 g499_reg ( .D(n6273), .CK(clk), .RN(n8025), .SN(1'b1), .Q(n12926) );
  DFFSRX1 g691_reg ( .D(n6272), .CK(clk), .RN(n8025), .SN(1'b1), .Q(n12920), 
        .QN(n7244) );
  DFFSRX1 g667_reg ( .D(n6271), .CK(clk), .RN(n8024), .SN(1'b1), .Q(n12329), 
        .QN(n7814) );
  DFFSRX1 g671_reg ( .D(n6270), .CK(clk), .RN(n8024), .SN(1'b1), .Q(n12170), 
        .QN(n7696) );
  DFFSRX1 g676_reg ( .D(n6269), .CK(clk), .RN(n8024), .SN(1'b1), .Q(n12168), 
        .QN(n7525) );
  DFFSRX1 g681_reg ( .D(n6268), .CK(clk), .RN(n8023), .SN(1'b1), .Q(n12178) );
  DFFSRX1 g699_reg ( .D(n6267), .CK(clk), .RN(n8023), .SN(1'b1), .Q(n7454), 
        .QN(n12179) );
  DFFSRX1 g703_reg ( .D(n6266), .CK(clk), .RN(n8025), .SN(1'b1), .Q(n12490), 
        .QN(n7407) );
  DFFSRX1 g837_reg ( .D(n6265), .CK(clk), .RN(n8025), .SN(1'b1), .Q(n7296), 
        .QN(n12165) );
  DFFSRX1 g843_reg ( .D(n6264), .CK(clk), .RN(n8024), .SN(1'b1), .QN(n7464) );
  DFFSRX1 g847_reg ( .D(n6263), .CK(clk), .RN(n8025), .SN(1'b1), .Q(n12166), 
        .QN(n7219) );
  DFFSRX1 g812_reg ( .D(n6262), .CK(clk), .RN(n8024), .SN(1'b1), .Q(n12167), 
        .QN(n7680) );
  DFFSRX1 g817_reg ( .D(n6261), .CK(clk), .RN(n8024), .SN(1'b1), .Q(n7357), 
        .QN(n12163) );
  DFFSRX1 g832_reg ( .D(n6260), .CK(clk), .RN(n8024), .SN(1'b1), .Q(n7368), 
        .QN(n12160) );
  DFFSRX1 g822_reg ( .D(n6259), .CK(clk), .RN(n8024), .SN(1'b1), .Q(n12164), 
        .QN(n7461) );
  DFFSRX1 g827_reg ( .D(n6258), .CK(clk), .RN(n8024), .SN(1'b1), .Q(n12161) );
  DFFSRX1 g723_reg ( .D(n6257), .CK(clk), .RN(n8023), .SN(1'b1), .Q(n12162), 
        .QN(n7630) );
  DFFSRX1 g732_reg ( .D(n6256), .CK(clk), .RN(n8085), .SN(1'b1), .Q(n12159) );
  DFFSRX1 g758_reg ( .D(n6255), .CK(clk), .RN(n8084), .SN(1'b1), .Q(n12224), 
        .QN(n7619) );
  DFFSRX1 g763_reg ( .D(n6254), .CK(clk), .RN(n8084), .SN(1'b1), .Q(n12223), 
        .QN(n7719) );
  DFFSRX1 g767_reg ( .D(n6253), .CK(clk), .RN(n8084), .SN(1'b1), .Q(n12222), 
        .QN(n7720) );
  DFFSRX1 g772_reg ( .D(n6252), .CK(clk), .RN(n8084), .SN(1'b1), .Q(n12221), 
        .QN(n7721) );
  DFFSRX1 g776_reg ( .D(n6251), .CK(clk), .RN(n8084), .SN(1'b1), .Q(n12220), 
        .QN(n7722) );
  DFFSRX1 g781_reg ( .D(n6250), .CK(clk), .RN(n8084), .SN(1'b1), .Q(n12219), 
        .QN(n7723) );
  DFFSRX1 g785_reg ( .D(n6249), .CK(clk), .RN(n8084), .SN(1'b1), .Q(n12218), 
        .QN(n7724) );
  DFFSRX1 g790_reg ( .D(n6248), .CK(clk), .RN(n8084), .SN(1'b1), .Q(n12217), 
        .QN(n7725) );
  DFFSRX1 g794_reg ( .D(n6247), .CK(clk), .RN(n8084), .SN(1'b1), .Q(n12228) );
  DFFSRX1 g802_reg ( .D(g12184), .CK(clk), .RN(n8085), .SN(1'b1), .Q(g11678), 
        .QN(n671) );
  DFFSRX1 g542_reg ( .D(n6246), .CK(clk), .RN(n8012), .SN(1'b1), .Q(n12247), 
        .QN(n7754) );
  DFFSRX1 g546_reg ( .D(n6245), .CK(clk), .RN(n8012), .SN(1'b1), .Q(n12242), 
        .QN(n7755) );
  DFFSRX1 g550_reg ( .D(n6244), .CK(clk), .RN(n8011), .SN(1'b1), .Q(n12950), 
        .QN(n7756) );
  DFFSRX1 g136_reg ( .D(n6243), .CK(clk), .RN(n7988), .SN(1'b1), .Q(g21292), 
        .QN(g30329) );
  DFFSRX1 g142_reg ( .D(n6242), .CK(clk), .RN(n7988), .SN(1'b1), .Q(n12914), 
        .QN(n7681) );
  DFFSRX1 g146_reg ( .D(n6241), .CK(clk), .RN(n8083), .SN(1'b1), .Q(n12904) );
  DFFSRX1 g150_reg ( .D(n6240), .CK(clk), .RN(n8083), .SN(1'b1), .Q(n12899), 
        .QN(n7682) );
  DFFSRX1 g153_reg ( .D(n6239), .CK(clk), .RN(n8083), .SN(1'b1), .Q(n12898), 
        .QN(n7726) );
  DFFSRX1 g157_reg ( .D(n6238), .CK(clk), .RN(n8083), .SN(1'b1), .Q(n12894), 
        .QN(n7727) );
  DFFSRX1 g160_reg ( .D(n6237), .CK(clk), .RN(n8083), .SN(1'b1), .QN(n7316) );
  DFFSRX1 g301_reg ( .D(n6236), .CK(clk), .RN(n8083), .SN(1'b1), .Q(n12777), 
        .QN(n7343) );
  DFFSRX1 g305_reg ( .D(n6235), .CK(clk), .RN(n8082), .SN(1'b1), .Q(n13060), 
        .QN(n7207) );
  DFFSRX1 g311_reg ( .D(n6234), .CK(clk), .RN(n8082), .SN(1'b1), .Q(n13058), 
        .QN(n7224) );
  DFFSRX1 g316_reg ( .D(n6233), .CK(clk), .RN(n8082), .SN(1'b1), .Q(n12590) );
  DFFSRX1 g319_reg ( .D(n6232), .CK(clk), .RN(n8082), .SN(1'b1), .Q(n7502), 
        .QN(n12589) );
  DFFSRX1 g329_reg ( .D(n6231), .CK(clk), .RN(n8082), .SN(1'b1), .Q(n13057), 
        .QN(n7811) );
  DFFSRX1 g333_reg ( .D(n6230), .CK(clk), .RN(n8082), .SN(1'b1), .Q(n12585), 
        .QN(n7342) );
  DFFSRX1 g336_reg ( .D(n6229), .CK(clk), .RN(n8082), .SN(1'b1), .Q(n12588), 
        .QN(n7520) );
  DFFSRX1 g324_reg ( .D(n6228), .CK(clk), .RN(n8082), .SN(1'b1), .Q(n13059), 
        .QN(n7283) );
  DFFSRX1 g358_reg ( .D(n6227), .CK(clk), .RN(n8027), .SN(1'b1), .Q(n12934) );
  DFFSRX1 g376_reg ( .D(n6226), .CK(clk), .RN(n8026), .SN(1'b1), .Q(n12933), 
        .QN(n7512) );
  DFFSRX1 g385_reg ( .D(n6225), .CK(clk), .RN(n8026), .SN(1'b1), .Q(n12932), 
        .QN(n7420) );
  DFFSRX1 g370_reg ( .D(n6224), .CK(clk), .RN(n8026), .SN(1'b1), .Q(n12931), 
        .QN(n7536) );
  DFFSRX1 g437_reg ( .D(n6223), .CK(clk), .RN(n8023), .SN(1'b1), .Q(n12476), 
        .QN(n7728) );
  DFFSRX1 g441_reg ( .D(n6222), .CK(clk), .RN(n8022), .SN(1'b1), .Q(n12439) );
  DFFSRX1 g446_reg ( .D(n6221), .CK(clk), .RN(n8022), .SN(1'b1), .Q(n12850), 
        .QN(n7606) );
  DFFSRX1 g417_reg ( .D(n6220), .CK(clk), .RN(n8023), .SN(1'b1), .Q(n12477), 
        .QN(n7370) );
  DFFSRX1 g424_reg ( .D(n6219), .CK(clk), .RN(n8023), .SN(1'b1), .Q(n12475), 
        .QN(n7321) );
  DFFSRX1 g401_reg ( .D(n6218), .CK(clk), .RN(n8013), .SN(1'b1), .Q(n12491), 
        .QN(n7729) );
  DFFSRX1 g392_reg ( .D(n6217), .CK(clk), .RN(n8023), .SN(1'b1), .Q(n12488), 
        .QN(n7373) );
  DFFSRX1 g405_reg ( .D(n6216), .CK(clk), .RN(n8013), .SN(1'b1), .Q(n12851) );
  DFFSRX1 g182_reg ( .D(n6215), .CK(clk), .RN(n8026), .SN(1'b1), .Q(n12903) );
  DFFSRX1 g191_reg ( .D(n6214), .CK(clk), .RN(n8012), .SN(1'b1), .Q(n12828), 
        .QN(n7631) );
  DFFSRX1 g194_reg ( .D(n6213), .CK(clk), .RN(n8012), .SN(1'b1), .Q(g8358), 
        .QN(n7800) );
  DFFSRX1 g209_reg ( .D(n6212), .CK(clk), .RN(n8012), .SN(1'b1), .Q(n12892) );
  DFFSRX1 g218_reg ( .D(g8291), .CK(clk), .RN(n8011), .SN(1'b1), .QN(n12829)
         );
  DFFSRX1 g225_reg ( .D(n6211), .CK(clk), .RN(n8085), .SN(1'b1), .Q(n12940), 
        .QN(n7223) );
  DFFSRX1 g255_reg ( .D(n6210), .CK(clk), .RN(n8014), .SN(1'b1), .Q(n12935), 
        .QN(n7222) );
  DFFSRX1 g232_reg ( .D(n6209), .CK(clk), .RN(n8013), .SN(1'b1), .Q(n12937), 
        .QN(n7281) );
  DFFSRX1 g262_reg ( .D(n6208), .CK(clk), .RN(n8013), .SN(1'b1), .Q(n12938), 
        .QN(n7286) );
  DFFSRX1 g239_reg ( .D(n6207), .CK(clk), .RN(n8013), .SN(1'b1), .Q(n12939), 
        .QN(n7397) );
  DFFSRX1 g269_reg ( .D(n6206), .CK(clk), .RN(n8013), .SN(1'b1), .Q(n7205), 
        .QN(n12936) );
  DFFSRX1 g246_reg ( .D(n6205), .CK(clk), .RN(n8013), .SN(1'b1), .Q(n13066), 
        .QN(n7206) );
  DFFSRX1 g278_reg ( .D(n6204), .CK(clk), .RN(n8013), .SN(1'b1), .QN(n7538) );
  DFFSRX1 g283_reg ( .D(n6203), .CK(clk), .RN(n8013), .SN(1'b1), .Q(n12919) );
  DFFSRX1 g287_reg ( .D(n6202), .CK(clk), .RN(n8012), .SN(1'b1), .Q(n7503), 
        .QN(n12918) );
  DFFSRX1 g291_reg ( .D(n6201), .CK(clk), .RN(n8012), .SN(1'b1), .Q(n12917) );
  DFFSRX1 g294_reg ( .D(n6200), .CK(clk), .RN(n8012), .SN(1'b1), .Q(n12916), 
        .QN(n7614) );
  DFFSRX1 g298_reg ( .D(n6199), .CK(clk), .RN(n8012), .SN(1'b1), .Q(n12915), 
        .QN(n7613) );
  DFFSRX1 g411_reg ( .D(n6198), .CK(clk), .RN(n8023), .SN(1'b1), .Q(n12478), 
        .QN(n7575) );
  DFFSRX1 g452_reg ( .D(n6197), .CK(clk), .RN(n8013), .SN(1'b1), .Q(n12415) );
  DFFSRX1 g460_reg ( .D(n6196), .CK(clk), .RN(n8013), .SN(1'b1), .Q(n12414) );
  DFFSRX1 g475_reg ( .D(n6195), .CK(clk), .RN(n8013), .SN(1'b1), .Q(n12435) );
  DFFSRX1 g513_reg ( .D(n6194), .CK(clk), .RN(n8083), .SN(1'b1), .Q(n12905), 
        .QN(n7615) );
  DFFSRX1 g518_reg ( .D(n6193), .CK(clk), .RN(n8026), .SN(1'b1), .Q(n12927), 
        .QN(n7605) );
  DFFSRX1 g479_reg ( .D(n6192), .CK(clk), .RN(n8026), .SN(1'b1), .Q(n7460) );
  DFFSRX1 g528_reg ( .D(n6191), .CK(clk), .RN(n8026), .SN(1'b1), .Q(n12930), 
        .QN(n7284) );
  DFFSRX1 g482_reg ( .D(n6190), .CK(clk), .RN(n8026), .SN(1'b1), .Q(n7365), 
        .QN(n12928) );
  DFFSRX1 g490_reg ( .D(n6189), .CK(clk), .RN(n8026), .SN(1'b1), .Q(n12929), 
        .QN(n7462) );
  DFFSRX1 g534_reg ( .D(n6188), .CK(clk), .RN(n8011), .SN(1'b1), .Q(n12246), 
        .QN(n7757) );
  DFFSRX1 g74_reg ( .D(n6187), .CK(clk), .RN(n8027), .SN(1'b1), .Q(g29211), 
        .QN(n5433) );
  DFFSRX1 g106_reg ( .D(n6186), .CK(clk), .RN(n8027), .SN(1'b1), .Q(g21176), 
        .QN(n5431) );
  DFFSRX1 g341_reg ( .D(n6185), .CK(clk), .RN(n8027), .SN(1'b1), .QN(n7820) );
  DFFSRX1 g344_reg ( .D(n6184), .CK(clk), .RN(n8027), .SN(1'b1), .Q(g7540), 
        .QN(n12533) );
  DFFSRX1 g347_reg ( .D(g7540), .CK(clk), .RN(n8027), .SN(1'b1), .QN(n7661) );
  DFFSRX1 g351_reg ( .D(n6183), .CK(clk), .RN(n8027), .SN(1'b1), .Q(n12158) );
  DFFSRX1 g128_reg ( .D(n6182), .CK(clk), .RN(n7988), .SN(1'b1), .Q(g21245), 
        .QN(n7647) );
  DFFSRX1 g2799_reg ( .D(n6181), .CK(clk), .RN(n7997), .SN(1'b1), .Q(n7302), 
        .QN(n12697) );
  DFFSRX1 g2803_reg ( .D(n6180), .CK(clk), .RN(n7991), .SN(1'b1), .Q(n7381), 
        .QN(n13020) );
  DFFSRX1 g2807_reg ( .D(n6179), .CK(clk), .RN(n7993), .SN(1'b1), .Q(n7378), 
        .QN(n13018) );
  DFFSRX1 g2811_reg ( .D(n6178), .CK(clk), .RN(n7997), .SN(1'b1), .Q(n7305), 
        .QN(n12688) );
  DFFSRX1 g2815_reg ( .D(n6177), .CK(clk), .RN(n7997), .SN(1'b1), .Q(n7271), 
        .QN(n13021) );
  DFFSRX1 g2819_reg ( .D(n6176), .CK(clk), .RN(n7997), .SN(1'b1), .Q(n7218), 
        .QN(n13019) );
  DFFSRX1 g2587_reg ( .D(n6175), .CK(clk), .RN(n7996), .SN(1'b1), .Q(n12711), 
        .QN(n7487) );
  DFFSRX1 g2638_reg ( .D(n6174), .CK(clk), .RN(n8009), .SN(1'b1), .Q(n13023), 
        .QN(n7325) );
  DFFSRX1 g2652_reg ( .D(n6173), .CK(clk), .RN(n8009), .SN(1'b1), .Q(n7435), 
        .QN(n12706) );
  DFFSRX1 g2657_reg ( .D(n6172), .CK(clk), .RN(n8009), .SN(1'b1), .Q(n12705), 
        .QN(n7216) );
  DFFSRX1 g2661_reg ( .D(n6171), .CK(clk), .RN(n8008), .SN(1'b1), .Q(n12704), 
        .QN(n7586) );
  DFFSRX1 g2667_reg ( .D(n6170), .CK(clk), .RN(n7996), .SN(1'b1), .Q(n12703)
         );
  DFFSRX1 g2671_reg ( .D(n6169), .CK(clk), .RN(n8008), .SN(1'b1), .QN(n7238)
         );
  DFFSRX1 g2675_reg ( .D(n6168), .CK(clk), .RN(n8008), .SN(1'b1), .Q(n12702), 
        .QN(n7308) );
  DFFSRX1 g2681_reg ( .D(n6167), .CK(clk), .RN(n7995), .SN(1'b1), .QN(n7662)
         );
  DFFSRX1 g2685_reg ( .D(n6166), .CK(clk), .RN(n8008), .SN(1'b1), .QN(n7213)
         );
  DFFSRX1 g2715_reg ( .D(n6165), .CK(clk), .RN(n8008), .SN(1'b1), .Q(n13032), 
        .QN(n7320) );
  DFFSRX1 g2719_reg ( .D(n6164), .CK(clk), .RN(n8008), .SN(1'b1), .Q(n13033), 
        .QN(n7574) );
  DFFSRX1 g2724_reg ( .D(n6163), .CK(clk), .RN(n8008), .SN(1'b1), .Q(n13028), 
        .QN(n7492) );
  DFFSRX1 g2729_reg ( .D(n6162), .CK(clk), .RN(n8008), .SN(1'b1), .Q(n13027), 
        .QN(n7300) );
  DFFSRX1 g2735_reg ( .D(n6161), .CK(clk), .RN(n8008), .SN(1'b1), .Q(n13026), 
        .QN(n7688) );
  DFFSRX1 g2741_reg ( .D(n6160), .CK(clk), .RN(n8008), .SN(1'b1), .Q(n13031), 
        .QN(n7319) );
  DFFSRX1 g2748_reg ( .D(n6159), .CK(clk), .RN(n8008), .SN(1'b1), .Q(n13029)
         );
  DFFSRX1 g2756_reg ( .D(n6158), .CK(clk), .RN(n8008), .SN(1'b1), .Q(n13030)
         );
  DFFSRX1 g2193_reg ( .D(n6157), .CK(clk), .RN(n7989), .SN(1'b1), .Q(n12783), 
        .QN(n7730) );
  DFFSRX1 g2197_reg ( .D(n6156), .CK(clk), .RN(n7989), .SN(1'b1), .Q(n12791), 
        .QN(n7465) );
  DFFSRX1 g2208_reg ( .D(n6155), .CK(clk), .RN(n7991), .SN(1'b1), .Q(n12781), 
        .QN(n7488) );
  DFFSRX1 g2217_reg ( .D(n6154), .CK(clk), .RN(n7991), .SN(1'b1), .Q(n12780), 
        .QN(n7290) );
  DFFSRX1 g2227_reg ( .D(n6153), .CK(clk), .RN(n7989), .SN(1'b1), .Q(n12793), 
        .QN(n7497) );
  DFFSRX1 g2165_reg ( .D(n6152), .CK(clk), .RN(n8011), .SN(1'b1), .Q(n12789)
         );
  DFFSRX1 g2161_reg ( .D(n6151), .CK(clk), .RN(n7989), .SN(1'b1), .Q(n12790)
         );
  DFFSRX1 g2169_reg ( .D(n6150), .CK(clk), .RN(n7989), .SN(1'b1), .Q(n12787)
         );
  DFFSRX1 g2173_reg ( .D(n6149), .CK(clk), .RN(n7988), .SN(1'b1), .Q(n12785)
         );
  DFFSRX1 g2177_reg ( .D(n6148), .CK(clk), .RN(n7989), .SN(1'b1), .Q(n12786)
         );
  DFFSRX1 g2181_reg ( .D(n6147), .CK(clk), .RN(n7989), .SN(1'b1), .Q(n7447), 
        .QN(n12784) );
  DFFSRX1 g2185_reg ( .D(n6146), .CK(clk), .RN(n7988), .SN(1'b1), .Q(n12782), 
        .QN(n7457) );
  DFFSRX1 g2259_reg ( .D(n6145), .CK(clk), .RN(n8011), .SN(1'b1), .Q(n12773), 
        .QN(n7587) );
  DFFSRX1 g2265_reg ( .D(n6144), .CK(clk), .RN(n7989), .SN(1'b1), .Q(n12768)
         );
  DFFSRX1 g2269_reg ( .D(n6143), .CK(clk), .RN(n8011), .SN(1'b1), .Q(n12767), 
        .QN(n7763) );
  DFFSRX1 g2273_reg ( .D(n6142), .CK(clk), .RN(n8011), .SN(1'b1), .Q(n12766), 
        .QN(n7521) );
  DFFSRX1 g2279_reg ( .D(n6141), .CK(clk), .RN(n8011), .SN(1'b1), .Q(n12765)
         );
  DFFSRX1 g2283_reg ( .D(n6140), .CK(clk), .RN(n8010), .SN(1'b1), .QN(n7335)
         );
  DFFSRX1 g2287_reg ( .D(n6139), .CK(clk), .RN(n8010), .SN(1'b1), .Q(n12763), 
        .QN(n7400) );
  DFFSRX1 g2380_reg ( .D(n6138), .CK(clk), .RN(n8010), .SN(1'b1), .Q(n12760)
         );
  DFFSRX1 g2299_reg ( .D(n6137), .CK(clk), .RN(n7991), .SN(1'b1), .Q(n12761)
         );
  DFFSRX1 g2303_reg ( .D(n6136), .CK(clk), .RN(n7991), .SN(1'b1), .Q(n12759)
         );
  DFFSRX1 g2315_reg ( .D(n6135), .CK(clk), .RN(n7993), .SN(1'b1), .Q(n7448), 
        .QN(n12756) );
  DFFSRX1 g2319_reg ( .D(n6134), .CK(clk), .RN(n7993), .SN(1'b1), .Q(n12753), 
        .QN(n7485) );
  DFFSRX1 g2327_reg ( .D(n6133), .CK(clk), .RN(n7993), .SN(1'b1), .Q(n12755), 
        .QN(n7731) );
  DFFSRX1 g2331_reg ( .D(n6132), .CK(clk), .RN(n7993), .SN(1'b1), .Q(n12762), 
        .QN(n7466) );
  DFFSRX1 g2295_reg ( .D(n6131), .CK(clk), .RN(n7991), .SN(1'b1), .Q(n7391) );
  DFFSRX1 g2342_reg ( .D(n6130), .CK(clk), .RN(n7993), .SN(1'b1), .Q(n12754), 
        .QN(n7550) );
  DFFSRX1 g2351_reg ( .D(n6129), .CK(clk), .RN(n7993), .SN(1'b1), .Q(n12752), 
        .QN(n7287) );
  DFFSRX1 g2361_reg ( .D(n6128), .CK(clk), .RN(n7993), .SN(1'b1), .Q(n12764)
         );
  DFFSRX1 g2307_reg ( .D(n6127), .CK(clk), .RN(n7991), .SN(1'b1), .Q(n12757)
         );
  DFFSRX1 g2311_reg ( .D(n6126), .CK(clk), .RN(n7991), .SN(1'b1), .Q(n12758)
         );
  DFFSRX1 g2370_reg ( .D(n6125), .CK(clk), .RN(n7991), .SN(1'b1), .Q(n13022), 
        .QN(n7594) );
  DFFSRX1 g2384_reg ( .D(n6124), .CK(clk), .RN(n7991), .SN(1'b1), .Q(n7436), 
        .QN(n12748) );
  DFFSRX1 g2389_reg ( .D(n6123), .CK(clk), .RN(n8010), .SN(1'b1), .Q(n12747), 
        .QN(n7351) );
  DFFSRX1 g2393_reg ( .D(n6122), .CK(clk), .RN(n8010), .SN(1'b1), .Q(n12746), 
        .QN(n7588) );
  DFFSRX1 g2399_reg ( .D(n6121), .CK(clk), .RN(n8010), .SN(1'b1), .Q(n12745)
         );
  DFFSRX1 g2403_reg ( .D(n6120), .CK(clk), .RN(n8010), .SN(1'b1), .QN(n7237)
         );
  DFFSRX1 g2407_reg ( .D(n6119), .CK(clk), .RN(n8010), .SN(1'b1), .Q(n12744), 
        .QN(n7309) );
  DFFSRX1 g2413_reg ( .D(n6118), .CK(clk), .RN(n7993), .SN(1'b1), .QN(n7663)
         );
  DFFSRX1 g2417_reg ( .D(n6117), .CK(clk), .RN(n8010), .SN(1'b1), .QN(n7212)
         );
  DFFSRX1 g2421_reg ( .D(n6116), .CK(clk), .RN(n8010), .SN(1'b1), .Q(n12742), 
        .QN(n7401) );
  DFFSRX1 g2514_reg ( .D(n6115), .CK(clk), .RN(n8009), .SN(1'b1), .Q(n12739)
         );
  DFFSRX1 g2433_reg ( .D(n6114), .CK(clk), .RN(n7998), .SN(1'b1), .Q(n12740)
         );
  DFFSRX1 g2437_reg ( .D(n6113), .CK(clk), .RN(n7995), .SN(1'b1), .Q(n12738)
         );
  DFFSRX1 g2449_reg ( .D(n6112), .CK(clk), .RN(n7995), .SN(1'b1), .Q(n7449), 
        .QN(n12735) );
  DFFSRX1 g2453_reg ( .D(n6111), .CK(clk), .RN(n7995), .SN(1'b1), .Q(n12732), 
        .QN(n7486) );
  DFFSRX1 g2461_reg ( .D(n6110), .CK(clk), .RN(n7998), .SN(1'b1), .Q(n12734), 
        .QN(n7735) );
  DFFSRX1 g2465_reg ( .D(n6109), .CK(clk), .RN(n7998), .SN(1'b1), .Q(n12741), 
        .QN(n7467) );
  DFFSRX1 g2429_reg ( .D(n6108), .CK(clk), .RN(n7998), .SN(1'b1), .Q(n7392) );
  DFFSRX1 g2476_reg ( .D(n6107), .CK(clk), .RN(n7995), .SN(1'b1), .Q(n12733), 
        .QN(n7552) );
  DFFSRX1 g2491_reg ( .D(n6106), .CK(clk), .RN(n7995), .SN(1'b1), .Q(n12729), 
        .QN(n7235) );
  DFFSRX1 g2485_reg ( .D(n6105), .CK(clk), .RN(n7995), .SN(1'b1), .Q(n12731), 
        .QN(n7288) );
  DFFSRX1 g2495_reg ( .D(n6104), .CK(clk), .RN(n7995), .SN(1'b1), .Q(n12743)
         );
  DFFSRX1 g2441_reg ( .D(n6103), .CK(clk), .RN(n7995), .SN(1'b1), .Q(n12736)
         );
  DFFSRX1 g2445_reg ( .D(n6102), .CK(clk), .RN(n7995), .SN(1'b1), .Q(n12737)
         );
  DFFSRX1 g2504_reg ( .D(n6101), .CK(clk), .RN(n7993), .SN(1'b1), .Q(n13024), 
        .QN(n7595) );
  DFFSRX1 g2518_reg ( .D(n6100), .CK(clk), .RN(n7993), .SN(1'b1), .Q(n7437), 
        .QN(n12727) );
  DFFSRX1 g2523_reg ( .D(n6099), .CK(clk), .RN(n8009), .SN(1'b1), .Q(n12726), 
        .QN(n7241) );
  DFFSRX1 g2527_reg ( .D(n6098), .CK(clk), .RN(n8009), .SN(1'b1), .Q(n12725), 
        .QN(n7589) );
  DFFSRX1 g2533_reg ( .D(n6097), .CK(clk), .RN(n8009), .SN(1'b1), .Q(n12724)
         );
  DFFSRX1 g2537_reg ( .D(n6096), .CK(clk), .RN(n8009), .SN(1'b1), .QN(n7648)
         );
  DFFSRX1 g2541_reg ( .D(n6095), .CK(clk), .RN(n8009), .SN(1'b1), .Q(n12723), 
        .QN(n7310) );
  DFFSRX1 g2547_reg ( .D(n6094), .CK(clk), .RN(n7995), .SN(1'b1), .QN(n7664)
         );
  DFFSRX1 g2551_reg ( .D(n6093), .CK(clk), .RN(n8009), .SN(1'b1), .QN(n7336)
         );
  DFFSRX1 g2555_reg ( .D(n6092), .CK(clk), .RN(n8009), .SN(1'b1), .Q(n12721), 
        .QN(n7402) );
  DFFSRX1 g2648_reg ( .D(n6091), .CK(clk), .RN(n7996), .SN(1'b1), .Q(n12718)
         );
  DFFSRX1 g2567_reg ( .D(n6090), .CK(clk), .RN(n7996), .SN(1'b1), .Q(n12719)
         );
  DFFSRX1 g2571_reg ( .D(n6089), .CK(clk), .RN(n7996), .SN(1'b1), .Q(n12717)
         );
  DFFSRX1 g2583_reg ( .D(n6088), .CK(clk), .RN(n7996), .SN(1'b1), .Q(n7450), 
        .QN(n12714) );
  DFFSRX1 g2579_reg ( .D(n6087), .CK(clk), .RN(n7996), .SN(1'b1), .Q(n12716)
         );
  DFFSRX1 g2575_reg ( .D(n6086), .CK(clk), .RN(n7995), .SN(1'b1), .Q(n12715)
         );
  DFFSRX1 g2595_reg ( .D(n6085), .CK(clk), .RN(n7996), .SN(1'b1), .Q(n12713), 
        .QN(n7736) );
  DFFSRX1 g2599_reg ( .D(n6084), .CK(clk), .RN(n7996), .SN(1'b1), .Q(n12720), 
        .QN(n7468) );
  DFFSRX1 g2563_reg ( .D(n6083), .CK(clk), .RN(n8009), .SN(1'b1), .Q(n7393) );
  DFFSRX1 g2610_reg ( .D(n6082), .CK(clk), .RN(n7997), .SN(1'b1), .Q(n12712), 
        .QN(n7553) );
  DFFSRX1 g2625_reg ( .D(n6081), .CK(clk), .RN(n7997), .SN(1'b1), .Q(n12708), 
        .QN(n7211) );
  DFFSRX1 g2619_reg ( .D(n6080), .CK(clk), .RN(n7997), .SN(1'b1), .Q(n12710), 
        .QN(n7289) );
  DFFSRX1 g2629_reg ( .D(n6079), .CK(clk), .RN(n7996), .SN(1'b1), .Q(n12722)
         );
  DFFSRX1 g2236_reg ( .D(n6078), .CK(clk), .RN(n8011), .SN(1'b1), .Q(n13025), 
        .QN(n7326) );
  DFFSRX1 g2759_reg ( .D(n6077), .CK(clk), .RN(n8007), .SN(1'b1), .QN(n7897)
         );
  DFFSRX1 g2787_reg ( .D(n6076), .CK(clk), .RN(n8005), .SN(1'b1), .Q(n13009), 
        .QN(n7531) );
  DFFSRX1 g2028_reg ( .D(n6075), .CK(clk), .RN(n7999), .SN(1'b1), .Q(n12804), 
        .QN(n7489) );
  DFFSRX1 g2036_reg ( .D(n6074), .CK(clk), .RN(n8005), .SN(1'b1), .Q(n12805), 
        .QN(n7687) );
  DFFSRX1 g2040_reg ( .D(n6073), .CK(clk), .RN(n8000), .SN(1'b1), .Q(n12818), 
        .QN(n7469) );
  DFFSRX1 g2047_reg ( .D(n6072), .CK(clk), .RN(n8000), .SN(1'b1), .Q(n12801), 
        .QN(n7346) );
  DFFSRX1 g2051_reg ( .D(n6071), .CK(clk), .RN(n7999), .SN(1'b1), .Q(n12803), 
        .QN(n7554) );
  DFFSRX1 g2066_reg ( .D(n6070), .CK(clk), .RN(n7999), .SN(1'b1), .Q(n12800), 
        .QN(n7209) );
  DFFSRX1 g2060_reg ( .D(n6069), .CK(clk), .RN(n7999), .SN(1'b1), .Q(n12802), 
        .QN(n7291) );
  DFFSRX1 g2070_reg ( .D(n6068), .CK(clk), .RN(n8000), .SN(1'b1), .Q(n12820)
         );
  DFFSRX1 g2008_reg ( .D(n6067), .CK(clk), .RN(n8000), .SN(1'b1), .Q(n12811)
         );
  DFFSRX1 g2004_reg ( .D(n6066), .CK(clk), .RN(n7999), .SN(1'b1), .Q(n7394) );
  DFFSRX1 g2012_reg ( .D(n6065), .CK(clk), .RN(n7999), .SN(1'b1), .Q(n12809)
         );
  DFFSRX1 g2024_reg ( .D(n6064), .CK(clk), .RN(n7999), .SN(1'b1), .Q(n7451), 
        .QN(n12806) );
  DFFSRX1 g2020_reg ( .D(n6063), .CK(clk), .RN(n7999), .SN(1'b1), .Q(n12808)
         );
  DFFSRX1 g2016_reg ( .D(n6062), .CK(clk), .RN(n7999), .SN(1'b1), .Q(n12807)
         );
  DFFSRX1 g2079_reg ( .D(n6061), .CK(clk), .RN(n8000), .SN(1'b1), .Q(n13013), 
        .QN(n7315) );
  DFFSRX1 g2791_reg ( .D(n6060), .CK(clk), .RN(n8001), .SN(1'b1), .Q(n7328), 
        .QN(n12699) );
  DFFSRX1 g2783_reg ( .D(n6059), .CK(clk), .RN(n8005), .SN(1'b1), .Q(n7414), 
        .QN(n13011) );
  DFFSRX1 g2775_reg ( .D(n6058), .CK(clk), .RN(n8005), .SN(1'b1), .Q(n7377), 
        .QN(n13008) );
  DFFSRX1 g2771_reg ( .D(n6057), .CK(clk), .RN(n8005), .SN(1'b1), .Q(n7297), 
        .QN(n13010) );
  DFFSRX1 g1677_reg ( .D(n6056), .CK(clk), .RN(n8005), .SN(1'b1), .Q(n13015), 
        .QN(n7617) );
  DFFSRX1 g1687_reg ( .D(n6055), .CK(clk), .RN(n8004), .SN(1'b1), .Q(n12886), 
        .QN(n7590) );
  DFFSRX1 g1604_reg ( .D(n6054), .CK(clk), .RN(n8004), .SN(1'b1), .Q(n12887)
         );
  DFFSRX1 g1608_reg ( .D(n6053), .CK(clk), .RN(n8004), .SN(1'b1), .Q(n12885)
         );
  DFFSRX1 g1620_reg ( .D(n6052), .CK(clk), .RN(n8004), .SN(1'b1), .Q(n7452), 
        .QN(n12882) );
  DFFSRX1 g1624_reg ( .D(n6051), .CK(clk), .RN(n8004), .SN(1'b1), .Q(n12880), 
        .QN(n7273) );
  DFFSRX1 g1632_reg ( .D(n6050), .CK(clk), .RN(n8004), .SN(1'b1), .Q(n12881), 
        .QN(n7733) );
  DFFSRX1 g2767_reg ( .D(n6049), .CK(clk), .RN(n8004), .SN(1'b1), .Q(n7304), 
        .QN(n12701) );
  DFFSRX1 g1636_reg ( .D(n6048), .CK(clk), .RN(n8004), .SN(1'b1), .Q(n12891), 
        .QN(n7421) );
  DFFSRX1 g1648_reg ( .D(n6047), .CK(clk), .RN(n8003), .SN(1'b1), .Q(n12879), 
        .QN(n7511) );
  DFFSRX1 g1657_reg ( .D(n6046), .CK(clk), .RN(n8003), .SN(1'b1), .Q(n12878), 
        .QN(n7404) );
  DFFSRX1 g1668_reg ( .D(n6045), .CK(clk), .RN(n8003), .SN(1'b1), .Q(n12890)
         );
  DFFSRX1 g1592_reg ( .D(n6044), .CK(clk), .RN(n8003), .SN(1'b1), .Q(n12889), 
        .QN(n7458) );
  DFFSRX1 g1616_reg ( .D(n6043), .CK(clk), .RN(n8004), .SN(1'b1), .Q(n12884)
         );
  DFFSRX1 g1612_reg ( .D(n6042), .CK(clk), .RN(n8004), .SN(1'b1), .Q(n12883)
         );
  DFFSRX1 g1600_reg ( .D(n6041), .CK(clk), .RN(n8004), .SN(1'b1), .Q(n12888)
         );
  DFFSRX1 g1691_reg ( .D(n6040), .CK(clk), .RN(n8003), .SN(1'b1), .Q(n12874), 
        .QN(n7314) );
  DFFSRX1 g1696_reg ( .D(n6039), .CK(clk), .RN(n8003), .SN(1'b1), .Q(n7602), 
        .QN(n12873) );
  DFFSRX1 g1700_reg ( .D(n6038), .CK(clk), .RN(n8003), .SN(1'b1), .Q(n12872), 
        .QN(n7591) );
  DFFSRX1 g1706_reg ( .D(n6037), .CK(clk), .RN(n8003), .SN(1'b1), .Q(n12871)
         );
  DFFSRX1 g1710_reg ( .D(n6036), .CK(clk), .RN(n8003), .SN(1'b1), .QN(n7337)
         );
  DFFSRX1 g1714_reg ( .D(n6035), .CK(clk), .RN(n8003), .SN(1'b1), .Q(n12870), 
        .QN(n7514) );
  DFFSRX1 g1720_reg ( .D(n6034), .CK(clk), .RN(n8003), .SN(1'b1), .Q(n12869)
         );
  DFFSRX1 g1724_reg ( .D(n6033), .CK(clk), .RN(n8002), .SN(1'b1), .QN(n7239)
         );
  DFFSRX1 g1728_reg ( .D(n6032), .CK(clk), .RN(n8002), .SN(1'b1), .Q(n12867), 
        .QN(n7405) );
  DFFSRX1 g1821_reg ( .D(n6031), .CK(clk), .RN(n8002), .SN(1'b1), .Q(n12864)
         );
  DFFSRX1 g1740_reg ( .D(n6030), .CK(clk), .RN(n8002), .SN(1'b1), .Q(n12865)
         );
  DFFSRX1 g1744_reg ( .D(n6029), .CK(clk), .RN(n8002), .SN(1'b1), .Q(n12863)
         );
  DFFSRX1 g1756_reg ( .D(n6028), .CK(clk), .RN(n8002), .SN(1'b1), .Q(n7453), 
        .QN(n12860) );
  DFFSRX1 g1760_reg ( .D(n6027), .CK(clk), .RN(n8002), .SN(1'b1), .Q(n12858), 
        .QN(n7490) );
  DFFSRX1 g1768_reg ( .D(n6026), .CK(clk), .RN(n8002), .SN(1'b1), .Q(n12859), 
        .QN(n7686) );
  DFFSRX1 g1772_reg ( .D(n6025), .CK(clk), .RN(n8001), .SN(1'b1), .Q(n12866), 
        .QN(n7470) );
  DFFSRX1 g1736_reg ( .D(n6024), .CK(clk), .RN(n8002), .SN(1'b1), .Q(n7395) );
  DFFSRX1 g1783_reg ( .D(n6023), .CK(clk), .RN(n8001), .SN(1'b1), .Q(n12857), 
        .QN(n7555) );
  DFFSRX1 g1792_reg ( .D(n6022), .CK(clk), .RN(n8001), .SN(1'b1), .Q(n12856), 
        .QN(n7292) );
  DFFSRX1 g1802_reg ( .D(n6021), .CK(clk), .RN(n8001), .SN(1'b1), .Q(n12868)
         );
  DFFSRX1 g1748_reg ( .D(n6020), .CK(clk), .RN(n8002), .SN(1'b1), .Q(n12861)
         );
  DFFSRX1 g1752_reg ( .D(n6019), .CK(clk), .RN(n8002), .SN(1'b1), .Q(n12862)
         );
  DFFSRX1 g1811_reg ( .D(n6018), .CK(clk), .RN(n8001), .SN(1'b1), .Q(n13012), 
        .QN(n7524) );
  DFFSRX1 g1825_reg ( .D(n6017), .CK(clk), .RN(n8001), .SN(1'b1), .Q(n12852), 
        .QN(n7522) );
  DFFSRX1 g1830_reg ( .D(n6016), .CK(clk), .RN(n8001), .SN(1'b1), .Q(n7603), 
        .QN(n12849) );
  DFFSRX1 g1834_reg ( .D(n6015), .CK(clk), .RN(n8001), .SN(1'b1), .Q(n12848), 
        .QN(n7592) );
  DFFSRX1 g1840_reg ( .D(n6014), .CK(clk), .RN(n8000), .SN(1'b1), .Q(n12847)
         );
  DFFSRX1 g1844_reg ( .D(n6013), .CK(clk), .RN(n8000), .SN(1'b1), .QN(n7214)
         );
  DFFSRX1 g1848_reg ( .D(n6012), .CK(clk), .RN(n8000), .SN(1'b1), .Q(n12846), 
        .QN(n7311) );
  DFFSRX1 g1854_reg ( .D(n6011), .CK(clk), .RN(n8000), .SN(1'b1), .QN(n7665)
         );
  DFFSRX1 g1858_reg ( .D(n6010), .CK(clk), .RN(n8000), .SN(1'b1), .Q(n12845), 
        .QN(n7764) );
  DFFSRX1 g1862_reg ( .D(n6009), .CK(clk), .RN(n8007), .SN(1'b1), .Q(n12843), 
        .QN(n7257) );
  DFFSRX1 g1955_reg ( .D(n6008), .CK(clk), .RN(n8006), .SN(1'b1), .Q(n12840)
         );
  DFFSRX1 g1874_reg ( .D(n6007), .CK(clk), .RN(n8007), .SN(1'b1), .Q(n12841)
         );
  DFFSRX1 g1878_reg ( .D(n6006), .CK(clk), .RN(n8007), .SN(1'b1), .Q(n12839)
         );
  DFFSRX1 g1890_reg ( .D(n6005), .CK(clk), .RN(n8006), .SN(1'b1), .Q(n7505), 
        .QN(n12836) );
  DFFSRX1 g1894_reg ( .D(n6004), .CK(clk), .RN(n8005), .SN(1'b1), .Q(n12834), 
        .QN(n7491) );
  DFFSRX1 g1902_reg ( .D(n6003), .CK(clk), .RN(n8007), .SN(1'b1), .Q(n12835), 
        .QN(n7732) );
  DFFSRX1 g1906_reg ( .D(n6002), .CK(clk), .RN(n8007), .SN(1'b1), .Q(n12842), 
        .QN(n7293) );
  DFFSRX1 g1870_reg ( .D(n6001), .CK(clk), .RN(n8007), .SN(1'b1), .Q(n7396) );
  DFFSRX1 g1917_reg ( .D(n6000), .CK(clk), .RN(n8007), .SN(1'b1), .Q(n12833), 
        .QN(n7556) );
  DFFSRX1 g1926_reg ( .D(n5999), .CK(clk), .RN(n8007), .SN(1'b1), .Q(n12832), 
        .QN(n7294) );
  DFFSRX1 g1936_reg ( .D(n5998), .CK(clk), .RN(n8007), .SN(1'b1), .Q(n12844), 
        .QN(n7510) );
  DFFSRX1 g1882_reg ( .D(n5997), .CK(clk), .RN(n8006), .SN(1'b1), .Q(n12837)
         );
  DFFSRX1 g1886_reg ( .D(n5996), .CK(clk), .RN(n8006), .SN(1'b1), .Q(n12838)
         );
  DFFSRX1 g2882_reg ( .D(n5995), .CK(clk), .RN(n8080), .SN(1'b1), .QN(n12666)
         );
  DFFSRX1 g2886_reg ( .D(n5994), .CK(clk), .RN(n8080), .SN(1'b1), .Q(n12662), 
        .QN(n7758) );
  DFFSRX1 g37_reg ( .D(n5993), .CK(clk), .RN(n8080), .SN(1'b1), .Q(g37), .QN(
        g23002) );
  DFFSRX1 g55_reg ( .D(n5992), .CK(clk), .RN(n8080), .SN(1'b1), .Q(n12536), 
        .QN(n7684) );
  DFFSRX1 g4531_reg ( .D(n5991), .CK(clk), .RN(n7987), .SN(1'b1), .QN(n7822)
         );
  DFFSRX1 g4534_reg ( .D(n5990), .CK(clk), .RN(n7985), .SN(1'b1), .Q(n12434)
         );
  DFFSRX1 g4423_reg ( .D(n5989), .CK(clk), .RN(n8079), .SN(1'b1), .Q(n12441), 
        .QN(n7734) );
  DFFSRX1 g4427_reg ( .D(n5988), .CK(clk), .RN(n7987), .SN(1'b1), .Q(n12675), 
        .QN(n7769) );
  DFFSRX1 g4434_reg ( .D(n5987), .CK(clk), .RN(n8077), .SN(1'b1), .Q(n12432), 
        .QN(n7632) );
  DFFSRX1 g4438_reg ( .D(n5986), .CK(clk), .RN(n8077), .SN(1'b1), .Q(n12430), 
        .QN(n7683) );
  DFFSRX1 g4449_reg ( .D(n5985), .CK(clk), .RN(n8077), .SN(1'b1), .Q(g7260), 
        .QN(n5304) );
  DFFSRX1 g4443_reg ( .D(n5984), .CK(clk), .RN(n8077), .SN(1'b1), .Q(n7600), 
        .QN(n12431) );
  DFFSRX1 g4452_reg ( .D(n5983), .CK(clk), .RN(n8076), .SN(1'b1), .Q(n12429)
         );
  DFFSRX1 g4459_reg ( .D(n5982), .CK(clk), .RN(n8076), .SN(1'b1), .Q(n12448), 
        .QN(n7633) );
  DFFSRX1 g4462_reg ( .D(n5981), .CK(clk), .RN(n8076), .SN(1'b1), .Q(n7228), 
        .QN(n12428) );
  DFFSRX1 g4467_reg ( .D(n5980), .CK(clk), .RN(n8076), .SN(1'b1), .Q(n12427), 
        .QN(n7530) );
  DFFSRX1 g4473_reg ( .D(n5979), .CK(clk), .RN(n8076), .SN(1'b1), .Q(n12449), 
        .QN(n7317) );
  DFFSRX1 g4369_reg ( .D(n5978), .CK(clk), .RN(n8076), .SN(1'b1), .Q(n12537), 
        .QN(n7767) );
  DFFSRX1 g4480_reg ( .D(n5977), .CK(clk), .RN(n7987), .SN(1'b1), .Q(n12423)
         );
  DFFSRX1 g4495_reg ( .D(n5976), .CK(clk), .RN(n7987), .SN(1'b1), .QN(n5293)
         );
  DFFSRX1 g4498_reg ( .D(n5975), .CK(clk), .RN(n7987), .SN(1'b1), .QN(n5292)
         );
  DFFSRX1 g4501_reg ( .D(n5974), .CK(clk), .RN(n7987), .SN(1'b1), .QN(n7881)
         );
  DFFSRX1 g4515_reg ( .D(n5973), .CK(clk), .RN(n8078), .SN(1'b1), .Q(n12447), 
        .QN(n7739) );
  DFFSRX1 g4375_reg ( .D(n5972), .CK(clk), .RN(n8078), .SN(1'b1), .Q(n7275), 
        .QN(n12815) );
  DFFSRX1 g4382_reg ( .D(n5971), .CK(clk), .RN(n8077), .SN(1'b1), .Q(n12437), 
        .QN(n7475) );
  DFFSRX1 g4388_reg ( .D(n5970), .CK(clk), .RN(n8077), .SN(1'b1), .Q(n12438), 
        .QN(n7616) );
  DFFSRX1 g4401_reg ( .D(n5969), .CK(clk), .RN(n8077), .SN(1'b1), .Q(n12436), 
        .QN(n7738) );
  DFFSRX1 g4405_reg ( .D(n5968), .CK(clk), .RN(n8077), .SN(1'b1), .Q(n12816), 
        .QN(n7760) );
  DFFSRX1 g4408_reg ( .D(n5967), .CK(clk), .RN(n8077), .SN(1'b1), .Q(g7243), 
        .QN(n5289) );
  DFFSRX1 g4411_reg ( .D(n5966), .CK(clk), .RN(n8077), .SN(1'b1), .Q(n12817), 
        .QN(n7344) );
  DFFSRX1 g4417_reg ( .D(n5965), .CK(clk), .RN(n8077), .SN(1'b1), .Q(n12813), 
        .QN(n7761) );
  DFFSRX1 g4392_reg ( .D(n5964), .CK(clk), .RN(n8077), .SN(1'b1), .Q(n12814), 
        .QN(n7263) );
  DFFSRX1 g4446_reg ( .D(n5963), .CK(clk), .RN(n8076), .SN(1'b1), .Q(g7245), 
        .QN(n5305) );
  DFFSRX1 g34_reg ( .D(n5962), .CK(clk), .RN(n8080), .SN(1'b1), .QN(n7352) );
  DFFSRX1 g4420_reg ( .D(n5961), .CK(clk), .RN(n7985), .SN(1'b1), .Q(n12676)
         );
  DFFSRX1 g4521_reg ( .D(n5960), .CK(clk), .RN(n8078), .SN(1'b1), .Q(n7456), 
        .QN(n12418) );
  DFFSRX1 g4527_reg ( .D(n5959), .CK(clk), .RN(n8078), .SN(1'b1), .Q(n12422), 
        .QN(n7597) );
  DFFSRX1 g4540_reg ( .D(n5958), .CK(clk), .RN(n8079), .SN(1'b1), .QN(n5281)
         );
  DFFSRX1 g4543_reg ( .D(n5957), .CK(clk), .RN(n8079), .SN(1'b1), .Q(n12409)
         );
  DFFSRX1 g4546_reg ( .D(n5956), .CK(clk), .RN(n8079), .SN(1'b1), .QN(n7877)
         );
  DFFSRX1 g4564_reg ( .D(n5955), .CK(clk), .RN(n7985), .SN(1'b1), .Q(n12410)
         );
  DFFSRX1 g4567_reg ( .D(n5954), .CK(clk), .RN(n8079), .SN(1'b1), .Q(n12408), 
        .QN(n7830) );
  DFFSRX1 g1945_reg ( .D(n5953), .CK(clk), .RN(n8006), .SN(1'b1), .Q(n13014), 
        .QN(n7324) );
  DFFSRX1 g1959_reg ( .D(n5952), .CK(clk), .RN(n8006), .SN(1'b1), .Q(n12825), 
        .QN(n7523) );
  DFFSRX1 g1964_reg ( .D(n5951), .CK(clk), .RN(n8006), .SN(1'b1), .Q(n7604), 
        .QN(n12824) );
  DFFSRX1 g1968_reg ( .D(n5950), .CK(clk), .RN(n8006), .SN(1'b1), .Q(n12823), 
        .QN(n7593) );
  DFFSRX1 g1974_reg ( .D(n5949), .CK(clk), .RN(n8006), .SN(1'b1), .Q(n12822)
         );
  DFFSRX1 g1978_reg ( .D(n5948), .CK(clk), .RN(n8006), .SN(1'b1), .QN(n7649)
         );
  DFFSRX1 g1982_reg ( .D(n5947), .CK(clk), .RN(n8006), .SN(1'b1), .Q(n12821), 
        .QN(n7312) );
  DFFSRX1 g1988_reg ( .D(n5946), .CK(clk), .RN(n8005), .SN(1'b1), .QN(n7666)
         );
  DFFSRX1 g1992_reg ( .D(n5945), .CK(clk), .RN(n8005), .SN(1'b1), .QN(n7338)
         );
  DFFSRX1 g2779_reg ( .D(n5944), .CK(clk), .RN(n8001), .SN(1'b1), .Q(n7303), 
        .QN(n12700) );
  DFFSRX1 g2795_reg ( .D(n5943), .CK(clk), .RN(n8005), .SN(1'b1), .Q(n12698)
         );
  DFFSRX1 g2823_reg ( .D(n5942), .CK(clk), .RN(n7998), .SN(1'b1), .Q(n7329), 
        .QN(n12687) );
  DFFSRX1 g2827_reg ( .D(n5941), .CK(clk), .RN(n7997), .SN(1'b1), .Q(n7306), 
        .QN(n12686) );
  DFFSRX1 g2831_reg ( .D(n5940), .CK(clk), .RN(n7997), .SN(1'b1), .Q(n13007), 
        .QN(g30331) );
  DFFSRX1 g2834_reg ( .D(n5939), .CK(clk), .RN(n7997), .SN(1'b1), .Q(g2834), 
        .QN(g23652) );
  DFFSRX1 g739_reg ( .D(n5938), .CK(clk), .RN(n8084), .SN(1'b1), .Q(n12227), 
        .QN(n7695) );
  DFFSRX1 g744_reg ( .D(n5937), .CK(clk), .RN(n8084), .SN(1'b1), .Q(n12226), 
        .QN(n7737) );
  DFFSRX1 g749_reg ( .D(n5936), .CK(clk), .RN(n8084), .SN(1'b1), .Q(n12225), 
        .QN(n7639) );
  DFFSRX1 g753_reg ( .D(n5935), .CK(clk), .RN(n8085), .SN(1'b1), .Q(n7385), 
        .QN(n12922) );
  DFFSRX1 g645_reg ( .D(n5934), .CK(clk), .RN(n8083), .SN(1'b1), .Q(n12186) );
  DFFSRX1 g650_reg ( .D(n5933), .CK(clk), .RN(n8023), .SN(1'b1), .Q(n12177) );
  DFFSRX1 g655_reg ( .D(n5932), .CK(clk), .RN(n8023), .SN(1'b1), .Q(n12921), 
        .QN(n7463) );
  DFFSRX1 g661_reg ( .D(n5931), .CK(clk), .RN(n8024), .SN(1'b1), .Q(n12171), 
        .QN(n7535) );
  DFFSRX1 g714_reg ( .D(n5930), .CK(clk), .RN(n8024), .SN(1'b1), .QN(n7540) );
  DFFSRX1 g718_reg ( .D(n5929), .CK(clk), .RN(n8024), .SN(1'b1), .Q(n7251), 
        .QN(n12923) );
  DFFSRX1 g6661_reg ( .D(n5928), .CK(clk), .RN(n8034), .SN(1'b1), .Q(g17688), 
        .QN(n5672) );
  DFFSRX1 g6668_reg ( .D(g17688), .CK(clk), .RN(n8033), .SN(1'b1), .Q(g17722), 
        .QN(n7805) );
  DFFSRX1 g6675_reg ( .D(n5927), .CK(clk), .RN(n8033), .SN(1'b1), .Q(g14828)
         );
  DFFSRX1 g6704_reg ( .D(n5926), .CK(clk), .RN(n8033), .SN(1'b1), .Q(g17778), 
        .QN(n5671) );
  DFFSRX1 g6723_reg ( .D(n5925), .CK(clk), .RN(n8032), .SN(1'b1), .Q(n12294), 
        .QN(n7818) );
  DFFSRX1 g6727_reg ( .D(n5924), .CK(clk), .RN(n8033), .SN(1'b1), .Q(n12298), 
        .QN(n7424) );
  DFFSRX1 g6490_reg ( .D(n5923), .CK(clk), .RN(n8033), .SN(1'b1), .Q(g9817), 
        .QN(n3812) );
  DFFSRX1 g6486_reg ( .D(n5922), .CK(clk), .RN(n8033), .SN(1'b1), .Q(g9743), 
        .QN(n7986) );
  DFFSRX1 g6732_reg ( .D(n5921), .CK(clk), .RN(n8032), .SN(1'b1), .QN(n7667)
         );
  DFFSRX1 g6736_reg ( .D(n5920), .CK(clk), .RN(n8032), .SN(1'b1), .Q(n12303)
         );
  DFFSRX1 g6741_reg ( .D(n5919), .CK(clk), .RN(n8032), .SN(1'b1), .Q(n7248), 
        .QN(n12304) );
  DFFSRX1 g6719_reg ( .D(n5918), .CK(clk), .RN(n8032), .SN(1'b1), .Q(g17764)
         );
  INVX1 U6314 ( .A(n7947), .Y(n7936) );
  INVX1 U6315 ( .A(n7948), .Y(n7938) );
  INVX1 U6316 ( .A(n7954), .Y(n7937) );
  INVX1 U6317 ( .A(n7950), .Y(n7935) );
  INVX1 U6318 ( .A(n7947), .Y(n7943) );
  INVX1 U6319 ( .A(n7948), .Y(n7942) );
  INVX1 U6320 ( .A(n7949), .Y(n7941) );
  INVX1 U6321 ( .A(n7954), .Y(n7940) );
  INVX1 U6322 ( .A(n7947), .Y(n7927) );
  INVX1 U6323 ( .A(n7953), .Y(n7926) );
  INVX1 U6324 ( .A(n7954), .Y(n7925) );
  INVX1 U6325 ( .A(n7952), .Y(n7924) );
  INVX1 U6326 ( .A(n7948), .Y(n7934) );
  INVX1 U6327 ( .A(n7947), .Y(n7932) );
  INVX1 U6328 ( .A(n7951), .Y(n7929) );
  INVX1 U6329 ( .A(n7947), .Y(n7931) );
  INVX1 U6330 ( .A(n7952), .Y(n7928) );
  INVX1 U6331 ( .A(n7946), .Y(n7930) );
  INVX1 U6332 ( .A(n7952), .Y(n7939) );
  INVX1 U6333 ( .A(n7947), .Y(n7944) );
  INVX1 U6334 ( .A(n8086), .Y(n8077) );
  INVX1 U6335 ( .A(n8103), .Y(n7995) );
  INVX1 U6336 ( .A(n8100), .Y(n8008) );
  INVX1 U6337 ( .A(n8099), .Y(n8009) );
  INVX1 U6338 ( .A(n8098), .Y(n8013) );
  INVX1 U6339 ( .A(n8089), .Y(n8084) );
  INVX1 U6340 ( .A(n8094), .Y(n8024) );
  INVX1 U6341 ( .A(n8097), .Y(n8015) );
  INVX1 U6342 ( .A(n8097), .Y(n8016) );
  INVX1 U6343 ( .A(n8091), .Y(n8046) );
  INVX1 U6344 ( .A(n8091), .Y(n8047) );
  INVX1 U6345 ( .A(n8089), .Y(n8054) );
  INVX1 U6346 ( .A(n8090), .Y(n8053) );
  INVX1 U6347 ( .A(n8087), .Y(n8073) );
  INVX1 U6348 ( .A(n8092), .Y(n8035) );
  INVX1 U6349 ( .A(n8088), .Y(n8061) );
  INVX1 U6350 ( .A(n8090), .Y(n8051) );
  INVX1 U6351 ( .A(n8088), .Y(n8062) );
  INVX1 U6352 ( .A(n8093), .Y(n8050) );
  INVX1 U6353 ( .A(n8094), .Y(n8041) );
  INVX1 U6354 ( .A(n8086), .Y(n8075) );
  INVX1 U6355 ( .A(n8092), .Y(n8049) );
  INVX1 U6356 ( .A(n8089), .Y(n8056) );
  INVX1 U6357 ( .A(n8089), .Y(n8055) );
  INVX1 U6358 ( .A(n8087), .Y(n8082) );
  INVX1 U6359 ( .A(n8102), .Y(n7999) );
  INVX1 U6360 ( .A(n8096), .Y(n8019) );
  INVX1 U6361 ( .A(n8096), .Y(n8020) );
  INVX1 U6362 ( .A(n8092), .Y(n8033) );
  INVX1 U6363 ( .A(n8086), .Y(n8076) );
  INVX1 U6364 ( .A(n8100), .Y(n8006) );
  INVX1 U6365 ( .A(n8101), .Y(n8001) );
  INVX1 U6366 ( .A(n8100), .Y(n8002) );
  INVX1 U6367 ( .A(n8101), .Y(n8003) );
  INVX1 U6368 ( .A(n8101), .Y(n8004) );
  INVX1 U6369 ( .A(n8101), .Y(n8005) );
  INVX1 U6370 ( .A(n8100), .Y(n8007) );
  INVX1 U6371 ( .A(n8103), .Y(n7996) );
  INVX1 U6372 ( .A(n8102), .Y(n7998) );
  INVX1 U6373 ( .A(n8103), .Y(n7993) );
  INVX1 U6374 ( .A(n8099), .Y(n8010) );
  INVX1 U6375 ( .A(n8102), .Y(n7991) );
  INVX1 U6376 ( .A(n8102), .Y(n7997) );
  INVX1 U6377 ( .A(n8099), .Y(n8011) );
  INVX1 U6378 ( .A(n8098), .Y(n8012) );
  INVX1 U6379 ( .A(n8095), .Y(n8023) );
  INVX1 U6380 ( .A(n8093), .Y(n8027) );
  INVX1 U6381 ( .A(n8093), .Y(n8083) );
  INVX1 U6382 ( .A(n8097), .Y(n8017) );
  INVX1 U6383 ( .A(n8098), .Y(n8014) );
  INVX1 U6384 ( .A(n8096), .Y(n8018) );
  INVX1 U6385 ( .A(n8095), .Y(n8022) );
  INVX1 U6386 ( .A(n8095), .Y(n8021) );
  INVX1 U6387 ( .A(n8094), .Y(n8026) );
  INVX1 U6388 ( .A(n8094), .Y(n8025) );
  INVX1 U6389 ( .A(n8100), .Y(n8038) );
  INVX1 U6390 ( .A(n8090), .Y(n8052) );
  INVX1 U6391 ( .A(rst), .Y(n8030) );
  INVX1 U6392 ( .A(n8088), .Y(n8070) );
  INVX1 U6393 ( .A(n8091), .Y(n8045) );
  INVX1 U6394 ( .A(n8097), .Y(n8044) );
  INVX1 U6395 ( .A(rst), .Y(n8071) );
  INVX1 U6396 ( .A(n8090), .Y(n8040) );
  INVX1 U6397 ( .A(n8087), .Y(n8072) );
  INVX1 U6398 ( .A(n8093), .Y(n8028) );
  INVX1 U6399 ( .A(n8087), .Y(n8074) );
  INVX1 U6400 ( .A(n8093), .Y(n8029) );
  INVX1 U6401 ( .A(n8092), .Y(n8034) );
  INVX1 U6402 ( .A(n8103), .Y(n8036) );
  INVX1 U6403 ( .A(n8089), .Y(n8031) );
  INVX1 U6404 ( .A(n8094), .Y(n8057) );
  INVX1 U6405 ( .A(n8090), .Y(n8059) );
  INVX1 U6406 ( .A(n8088), .Y(n8060) );
  INVX1 U6407 ( .A(n8089), .Y(n8063) );
  INVX1 U6408 ( .A(n8086), .Y(n8064) );
  INVX1 U6409 ( .A(n8095), .Y(n8066) );
  INVX1 U6410 ( .A(n8101), .Y(n8065) );
  INVX1 U6411 ( .A(n8088), .Y(n8048) );
  INVX1 U6412 ( .A(n8091), .Y(n8039) );
  INVX1 U6413 ( .A(n8098), .Y(n8042) );
  INVX1 U6414 ( .A(n8096), .Y(n8043) );
  INVX1 U6415 ( .A(n8098), .Y(n8078) );
  INVX1 U6416 ( .A(n8102), .Y(n8037) );
  INVX1 U6417 ( .A(n8086), .Y(n8032) );
  INVX1 U6418 ( .A(n8099), .Y(n8067) );
  INVX1 U6419 ( .A(n8101), .Y(n8068) );
  INVX1 U6420 ( .A(n8087), .Y(n8069) );
  INVX1 U6421 ( .A(n8092), .Y(n8081) );
  INVX1 U6422 ( .A(n8096), .Y(n8079) );
  INVX1 U6423 ( .A(n8091), .Y(n8058) );
  INVX1 U6424 ( .A(n8099), .Y(n7988) );
  INVX1 U6425 ( .A(n8095), .Y(n8080) );
  INVX1 U6426 ( .A(n8097), .Y(n7989) );
  INVX1 U6427 ( .A(n8103), .Y(n8000) );
  INVX1 U6428 ( .A(n8086), .Y(n8085) );
  INVX1 U6429 ( .A(n7949), .Y(n7923) );
  INVX1 U6430 ( .A(n7946), .Y(n7945) );
  INVX1 U6431 ( .A(rst), .Y(n7987) );
  INVX1 U6432 ( .A(rst), .Y(n7985) );
  INVX1 U6433 ( .A(n7951), .Y(n7922) );
  INVX1 U6434 ( .A(n7916), .Y(n7874) );
  INVX1 U6435 ( .A(n7916), .Y(n7875) );
  INVX1 U6436 ( .A(n7917), .Y(n7876) );
  INVX1 U6437 ( .A(n7917), .Y(n7878) );
  INVX1 U6438 ( .A(n7916), .Y(n7879) );
  INVX1 U6439 ( .A(n7917), .Y(n7880) );
  INVX1 U6440 ( .A(n7916), .Y(n7882) );
  INVX1 U6441 ( .A(n7916), .Y(n7883) );
  INVX1 U6442 ( .A(n7916), .Y(n7884) );
  INVX1 U6443 ( .A(n7917), .Y(n7885) );
  INVX1 U6444 ( .A(n7916), .Y(n7886) );
  INVX1 U6445 ( .A(n7917), .Y(n7887) );
  INVX1 U6446 ( .A(n7917), .Y(n7888) );
  INVX1 U6447 ( .A(n7917), .Y(n7889) );
  INVX1 U6448 ( .A(n7917), .Y(n7890) );
  INVX1 U6449 ( .A(n7917), .Y(n7891) );
  INVX1 U6450 ( .A(n7917), .Y(n7892) );
  INVX1 U6451 ( .A(n7916), .Y(n7893) );
  INVX1 U6452 ( .A(n7916), .Y(n7894) );
  INVX1 U6453 ( .A(n7916), .Y(n7895) );
  INVX1 U6454 ( .A(n7917), .Y(n7896) );
  INVX1 U6455 ( .A(n7916), .Y(n7898) );
  INVX1 U6456 ( .A(n7916), .Y(n7899) );
  INVX1 U6457 ( .A(n7916), .Y(n7900) );
  INVX1 U6458 ( .A(n7917), .Y(n7901) );
  INVX1 U6459 ( .A(n7916), .Y(n7902) );
  INVX1 U6460 ( .A(n7916), .Y(n7903) );
  INVX1 U6461 ( .A(n7917), .Y(n7904) );
  INVX1 U6462 ( .A(n7916), .Y(n7905) );
  INVX1 U6463 ( .A(n7917), .Y(n7906) );
  INVX1 U6464 ( .A(n7916), .Y(n7907) );
  INVX1 U6465 ( .A(n7917), .Y(n7873) );
  INVX1 U6466 ( .A(n7917), .Y(n7908) );
  INVX1 U6467 ( .A(n7917), .Y(n7909) );
  INVX1 U6468 ( .A(n7916), .Y(n7914) );
  INVX1 U6469 ( .A(n7917), .Y(n7915) );
  INVX1 U6470 ( .A(n7917), .Y(n7913) );
  INVX1 U6471 ( .A(n7917), .Y(n7910) );
  INVX1 U6472 ( .A(n7871), .Y(n7860) );
  INVX1 U6473 ( .A(n7872), .Y(n7865) );
  INVX1 U6474 ( .A(n7872), .Y(n7866) );
  INVX1 U6475 ( .A(n7871), .Y(n7867) );
  INVX1 U6476 ( .A(n7871), .Y(n7868) );
  INVX1 U6477 ( .A(n7872), .Y(n7869) );
  INVX1 U6478 ( .A(n7871), .Y(n7870) );
  INVX1 U6479 ( .A(n7871), .Y(n7855) );
  INVX1 U6480 ( .A(n7872), .Y(n7857) );
  INVX1 U6481 ( .A(n7872), .Y(n7859) );
  INVX1 U6482 ( .A(n7872), .Y(n7856) );
  INVX1 U6483 ( .A(n7872), .Y(n7858) );
  INVX1 U6484 ( .A(n7872), .Y(n7854) );
  INVX1 U6485 ( .A(n7872), .Y(n7845) );
  INVX1 U6486 ( .A(n7871), .Y(n7852) );
  INVX1 U6487 ( .A(n7871), .Y(n7853) );
  INVX1 U6488 ( .A(n7872), .Y(n7846) );
  INVX1 U6489 ( .A(n7871), .Y(n7848) );
  INVX1 U6490 ( .A(n7871), .Y(n7849) );
  INVX1 U6491 ( .A(n7871), .Y(n7851) );
  INVX1 U6492 ( .A(n7871), .Y(n7850) );
  INVX1 U6493 ( .A(n7871), .Y(n7847) );
  INVX1 U6494 ( .A(n8114), .Y(n7976) );
  INVX1 U6495 ( .A(n8114), .Y(n7978) );
  INVX1 U6496 ( .A(n8114), .Y(n7963) );
  INVX1 U6497 ( .A(n8114), .Y(n7970) );
  INVX1 U6498 ( .A(n8114), .Y(n7971) );
  INVX1 U6499 ( .A(n8114), .Y(n7972) );
  INVX1 U6500 ( .A(n8114), .Y(n7974) );
  INVX1 U6501 ( .A(n8114), .Y(n7979) );
  INVX1 U6502 ( .A(n8114), .Y(n7969) );
  INVX1 U6503 ( .A(n8114), .Y(n7968) );
  INVX1 U6504 ( .A(n8114), .Y(n7980) );
  INVX1 U6505 ( .A(n8114), .Y(n7981) );
  INVX1 U6506 ( .A(n8114), .Y(n7982) );
  INVX1 U6507 ( .A(n8114), .Y(n7983) );
  INVX1 U6508 ( .A(n8114), .Y(n7962) );
  INVX1 U6509 ( .A(n8114), .Y(n7964) );
  INVX1 U6510 ( .A(n8114), .Y(n7965) );
  INVX1 U6511 ( .A(n8114), .Y(n7966) );
  INVX1 U6512 ( .A(n8114), .Y(n7967) );
  INVX1 U6513 ( .A(n8114), .Y(n7977) );
  INVX1 U6514 ( .A(n8114), .Y(n7961) );
  INVX1 U6515 ( .A(n8114), .Y(n7956) );
  INVX1 U6516 ( .A(n8114), .Y(n7959) );
  INVX1 U6517 ( .A(n8114), .Y(n7957) );
  INVX1 U6518 ( .A(n8114), .Y(n7958) );
  INVX1 U6519 ( .A(n8114), .Y(n7960) );
  INVX1 U6520 ( .A(n8114), .Y(n7955) );
  INVX1 U6521 ( .A(n8114), .Y(n7946) );
  INVX1 U6522 ( .A(n8114), .Y(n7952) );
  INVX1 U6523 ( .A(n8114), .Y(n7947) );
  INVX1 U6524 ( .A(n8114), .Y(n7948) );
  INVX1 U6525 ( .A(n8114), .Y(n7949) );
  INVX1 U6526 ( .A(n8114), .Y(n7950) );
  INVX1 U6527 ( .A(n8114), .Y(n7953) );
  INVX1 U6528 ( .A(n8114), .Y(n7954) );
  INVX1 U6529 ( .A(n8114), .Y(n7951) );
  INVX1 U6530 ( .A(n5917), .Y(n8089) );
  INVX1 U6531 ( .A(n5917), .Y(n8086) );
  INVX1 U6532 ( .A(n5917), .Y(n8101) );
  INVX1 U6533 ( .A(n5917), .Y(n8100) );
  INVX1 U6534 ( .A(n5917), .Y(n8103) );
  INVX1 U6535 ( .A(n5917), .Y(n8102) );
  INVX1 U6536 ( .A(n5917), .Y(n8099) );
  INVX1 U6537 ( .A(n5917), .Y(n8097) );
  INVX1 U6538 ( .A(n5917), .Y(n8098) );
  INVX1 U6539 ( .A(n5917), .Y(n8096) );
  INVX1 U6540 ( .A(n5917), .Y(n8095) );
  INVX1 U6541 ( .A(n5917), .Y(n8094) );
  INVX1 U6542 ( .A(n5917), .Y(n8090) );
  INVX1 U6543 ( .A(n5917), .Y(n8091) );
  INVX1 U6544 ( .A(n5917), .Y(n8087) );
  INVX1 U6545 ( .A(n5917), .Y(n8093) );
  INVX1 U6546 ( .A(n5917), .Y(n8092) );
  INVX1 U6547 ( .A(n5917), .Y(n8088) );
  INVX1 U6548 ( .A(n8108), .Y(n7919) );
  INVX1 U6549 ( .A(n8108), .Y(n7918) );
  INVX1 U6550 ( .A(n8108), .Y(n7920) );
  INVX1 U6551 ( .A(n8108), .Y(n7917) );
  INVX1 U6552 ( .A(n8108), .Y(n7916) );
  INVX1 U6553 ( .A(n8108), .Y(n7921) );
  INVX1 U6554 ( .A(n8104), .Y(n7872) );
  INVX1 U6555 ( .A(n8104), .Y(n7871) );
  OAI21X1 U6556 ( .A0(n7766), .A1(n7859), .B0(n8105), .Y(n7202) );
  MX2X1 U6557 ( .A(n8106), .B(n8107), .S0(n7623), .Y(n8105) );
  OR2X1 U6558 ( .A(n7969), .B(n5212), .Y(n8107) );
  AOI21X1 U6559 ( .A0(n5212), .A1(n7855), .B0(n8108), .Y(n8106) );
  MX2X1 U6560 ( .A(n8109), .B(test_se), .S0(n12934), .Y(n7201) );
  NOR2X1 U6561 ( .A(n7969), .B(g8719), .Y(n8109) );
  OAI21X1 U6562 ( .A0(n7921), .A1(n7420), .B0(n8110), .Y(n7200) );
  MX2X1 U6563 ( .A(n7800), .B(n8111), .S0(n7852), .Y(n8110) );
  OAI21X1 U6564 ( .A0(n5433), .A1(n7854), .B0(n8112), .Y(n7199) );
  AOI22X1 U6565 ( .A0(n8113), .A1(n7934), .B0(n12169), .B1(n8115), .Y(n8112)
         );
  OAI21X1 U6566 ( .A0(test_se), .A1(n8116), .B0(n7918), .Y(n8115) );
  MX2X1 U6567 ( .A(n12171), .B(g29212), .S0(n8116), .Y(n8113) );
  OAI21X1 U6568 ( .A0(n5870), .A1(n7854), .B0(n8117), .Y(n7198) );
  AOI22X1 U6569 ( .A0(n8108), .A1(n7460), .B0(n13066), .B1(n7931), .Y(n8117)
         );
  OAI21X1 U6570 ( .A0(n7854), .A1(n7462), .B0(n8118), .Y(n7197) );
  AOI22X1 U6571 ( .A0(n8108), .A1(g29215), .B0(n7928), .B1(n7205), .Y(n8118)
         );
  OAI21X1 U6572 ( .A0(n12829), .A1(n7854), .B0(n8119), .Y(n7196) );
  AOI22X1 U6573 ( .A0(n8120), .A1(n12914), .B0(n12777), .B1(n8108), .Y(n8119)
         );
  AND2X1 U6574 ( .A(n7928), .B(n8121), .Y(n8120) );
  OAI21X1 U6575 ( .A0(n7854), .A1(n7629), .B0(n8122), .Y(n7195) );
  NAND4X1 U6576 ( .A(n7911), .B(n699), .C(n8123), .D(n5266), .Y(n8122) );
  AOI21X1 U6577 ( .A0(n8124), .A1(n12944), .B0(n7969), .Y(n8123) );
  AOI21X1 U6578 ( .A0(n8125), .A1(n8126), .B0(n8127), .Y(n8124) );
  OAI21X1 U6579 ( .A0(n7855), .A1(n7628), .B0(n8128), .Y(n7194) );
  NAND4X1 U6580 ( .A(n7933), .B(n7912), .C(n8129), .D(n5246), .Y(n8128) );
  AOI21X1 U6581 ( .A0(n8130), .A1(n13049), .B0(n7969), .Y(n8129) );
  AOI21X1 U6582 ( .A0(n8131), .A1(n8132), .B0(n8133), .Y(n8130) );
  NAND2X1 U6583 ( .A(n7897), .B(n7969), .Y(n7193) );
  OAI21X1 U6584 ( .A0(n5239), .A1(n7854), .B0(n8134), .Y(n7192) );
  AOI21X1 U6585 ( .A0(n8108), .A1(n7353), .B0(n8135), .Y(n8134) );
  NOR2X1 U6586 ( .A(n8136), .B(n8137), .Y(n8135) );
  NAND4X1 U6587 ( .A(n12442), .B(n12443), .C(n12444), .D(n12445), .Y(n8137) );
  NAND4X1 U6588 ( .A(n12446), .B(n8138), .C(n8139), .D(n7412), .Y(n8136) );
  INVX1 U6589 ( .A(n8140), .Y(n8138) );
  OAI21X1 U6590 ( .A0(n5532), .A1(n7854), .B0(n8141), .Y(n7191) );
  AOI22X1 U6591 ( .A0(g37), .A1(n8108), .B0(n7928), .B1(g20652), .Y(n8141) );
  OAI21X1 U6592 ( .A0(n7855), .A1(n7767), .B0(n8142), .Y(n7190) );
  AOI21X1 U6593 ( .A0(n12538), .A1(n7891), .B0(n8143), .Y(n8142) );
  NOR2X1 U6594 ( .A(n8144), .B(n7969), .Y(n8143) );
  AOI21X1 U6595 ( .A0(n8145), .A1(n12453), .B0(n8146), .Y(n8144) );
  MX2X1 U6596 ( .A(n8147), .B(n8148), .S0(n7353), .Y(n8146) );
  NOR2X1 U6597 ( .A(n12452), .B(n12453), .Y(n8148) );
  NOR2X1 U6598 ( .A(n8149), .B(n7409), .Y(n8147) );
  AOI21X1 U6599 ( .A0(n8149), .A1(n12451), .B0(n8150), .Y(n8145) );
  INVX1 U6600 ( .A(n8151), .Y(n8149) );
  NAND3X1 U6601 ( .A(n12453), .B(n12452), .C(n8152), .Y(n8151) );
  MX2X1 U6602 ( .A(n8153), .B(n8154), .S0(n7364), .Y(n8152) );
  NAND2X1 U6603 ( .A(n12540), .B(n7375), .Y(n8154) );
  NAND2X1 U6604 ( .A(n7252), .B(n7739), .Y(n8153) );
  NAND2X1 U6605 ( .A(n7881), .B(n8155), .Y(n7189) );
  OAI21X1 U6606 ( .A0(n7928), .A1(n7739), .B0(n8156), .Y(n7188) );
  AOI22X1 U6607 ( .A0(n12417), .A1(n8157), .B0(n8158), .B1(g20049), .Y(n8156)
         );
  NAND2X1 U6608 ( .A(n8159), .B(n8160), .Y(n7187) );
  INVX1 U6609 ( .A(n8161), .Y(n8160) );
  MX2X1 U6610 ( .A(n12434), .B(n8162), .S0(n7853), .Y(n8161) );
  AOI21X1 U6611 ( .A0(n12424), .A1(n7893), .B0(n8163), .Y(n8159) );
  NAND2X1 U6612 ( .A(n8164), .B(n8165), .Y(n7186) );
  NAND2X1 U6613 ( .A(test_si), .B(test_se), .Y(n8165) );
  AOI22X1 U6614 ( .A0(n7928), .A1(n8166), .B0(n12812), .B1(n7883), .Y(n8164)
         );
  OAI21X1 U6615 ( .A0(n7855), .A1(n7344), .B0(n8167), .Y(n7185) );
  AOI22X1 U6616 ( .A0(n8168), .A1(n8169), .B0(n8170), .B1(n7275), .Y(n8167) );
  NAND2X1 U6617 ( .A(n8171), .B(n7969), .Y(n7184) );
  MX2X1 U6618 ( .A(n7758), .B(n7350), .S0(n7853), .Y(n8171) );
  OAI21X1 U6619 ( .A0(n7854), .A1(n7697), .B0(n8172), .Y(n7183) );
  AOI22X1 U6620 ( .A0(n12465), .A1(n7913), .B0(n7928), .B1(n7650), .Y(n8172)
         );
  OAI21X1 U6621 ( .A0(n5242), .A1(n7854), .B0(n8173), .Y(n7182) );
  AOI22X1 U6622 ( .A0(n8174), .A1(n7928), .B0(n7903), .B1(n7598), .Y(n8173) );
  MX2X1 U6623 ( .A(n7516), .B(n8175), .S0(n5240), .Y(n8174) );
  OAI21X1 U6624 ( .A0(n8176), .A1(n8177), .B0(n7516), .Y(n8175) );
  NAND3X1 U6625 ( .A(n7863), .B(n7862), .C(n7864), .Y(n8177) );
  NAND4X1 U6626 ( .A(n7861), .B(n5243), .C(n5242), .D(n5241), .Y(n8176) );
  OAI21X1 U6627 ( .A0(n5265), .A1(n7855), .B0(n8178), .Y(n7181) );
  AOI22X1 U6628 ( .A0(n7928), .A1(n8179), .B0(n13007), .B1(n7915), .Y(n8178)
         );
  OAI21X1 U6629 ( .A0(n5431), .A1(n7854), .B0(n8180), .Y(n7180) );
  AOI22X1 U6630 ( .A0(n7928), .A1(n8181), .B0(g2834), .B1(n7915), .Y(n8180) );
  NAND2X1 U6631 ( .A(n8182), .B(n7969), .Y(n7179) );
  MX2X1 U6632 ( .A(n7350), .B(n12666), .S0(n7852), .Y(n8182) );
  INVX1 U6633 ( .A(n8183), .Y(n7178) );
  AOI21X1 U6634 ( .A0(n7915), .A1(n12393), .B0(n8184), .Y(n8183) );
  MX2X1 U6635 ( .A(n12406), .B(n8185), .S0(n7852), .Y(n8184) );
  INVX1 U6636 ( .A(n8186), .Y(n7177) );
  AOI21X1 U6637 ( .A0(g20049), .A1(n7915), .B0(n8187), .Y(n8186) );
  MX2X1 U6638 ( .A(n12393), .B(n8188), .S0(n7854), .Y(n8187) );
  NAND2X1 U6639 ( .A(n7877), .B(n8155), .Y(n7176) );
  OAI21X1 U6640 ( .A0(n7855), .A1(n7830), .B0(n8189), .Y(n7175) );
  AOI22X1 U6641 ( .A0(n12407), .A1(n8190), .B0(n12406), .B1(n8158), .Y(n8189)
         );
  OAI21X1 U6642 ( .A0(test_se), .A1(n12425), .B0(n7918), .Y(n8190) );
  OAI21X1 U6643 ( .A0(n7855), .A1(n7757), .B0(n8191), .Y(n7174) );
  OAI21X1 U6644 ( .A0(n12892), .A1(n12245), .B0(n7922), .Y(n8191) );
  OAI21X1 U6645 ( .A0(n7856), .A1(n7768), .B0(n8192), .Y(n7173) );
  OAI21X1 U6646 ( .A0(n12650), .A1(n12639), .B0(n7922), .Y(n8192) );
  OAI21X1 U6647 ( .A0(n7855), .A1(n7769), .B0(n8193), .Y(n7172) );
  AOI21X1 U6648 ( .A0(n7928), .A1(n7600), .B0(n8194), .Y(n8193) );
  AOI21X1 U6649 ( .A0(n7921), .A1(n8195), .B0(n7632), .Y(n8194) );
  NAND3X1 U6650 ( .A(n12814), .B(n7856), .C(n8196), .Y(n8195) );
  OAI21X1 U6651 ( .A0(n7856), .A1(n7698), .B0(n8197), .Y(n7171) );
  AOI22X1 U6652 ( .A0(n8198), .A1(n8199), .B0(n12301), .B1(n8200), .Y(n8197)
         );
  OAI21X1 U6653 ( .A0(n7969), .A1(n8201), .B0(n8202), .Y(n8200) );
  AOI21X1 U6654 ( .A0(n8203), .A1(n8204), .B0(n8201), .Y(n8198) );
  MX2X1 U6655 ( .A(n8205), .B(n8206), .S0(n12529), .Y(n8204) );
  MX2X1 U6656 ( .A(n8207), .B(n8208), .S0(n12530), .Y(n8203) );
  OAI21X1 U6657 ( .A0(n7856), .A1(n7630), .B0(n8209), .Y(n7170) );
  AOI22X1 U6658 ( .A0(n12171), .A1(n8210), .B0(n8211), .B1(n12169), .Y(n8209)
         );
  OAI21X1 U6659 ( .A0(n7856), .A1(n7699), .B0(n8212), .Y(n7169) );
  AOI22X1 U6660 ( .A0(n8213), .A1(n8214), .B0(n12379), .B1(n8215), .Y(n8212)
         );
  AOI21X1 U6661 ( .A0(n7669), .A1(n8216), .B0(n7969), .Y(n8213) );
  OAI21X1 U6662 ( .A0(n8217), .A1(n8218), .B0(n8219), .Y(n8216) );
  MX2X1 U6663 ( .A(n8220), .B(n8221), .S0(n12376), .Y(n8218) );
  MX2X1 U6664 ( .A(n8222), .B(n8223), .S0(n7659), .Y(n8217) );
  NAND2X1 U6665 ( .A(n8224), .B(n8225), .Y(n7168) );
  MX2X1 U6666 ( .A(n8226), .B(n8227), .S0(n12909), .Y(n8225) );
  AOI21X1 U6667 ( .A0(n8228), .A1(n8229), .B0(test_se), .Y(n8227) );
  NAND2X1 U6668 ( .A(n8230), .B(n8228), .Y(n8226) );
  INVX1 U6669 ( .A(n8231), .Y(n8228) );
  AOI22X1 U6670 ( .A0(n8232), .A1(n8233), .B0(n12910), .B1(n7928), .Y(n8231)
         );
  AOI22X1 U6671 ( .A0(n8234), .A1(n12910), .B0(n12913), .B1(n7915), .Y(n8224)
         );
  NOR2X1 U6672 ( .A(n8233), .B(n7968), .Y(n8234) );
  NAND2X1 U6673 ( .A(n8235), .B(n8236), .Y(n7167) );
  MX2X1 U6674 ( .A(n8237), .B(n8238), .S0(n7367), .Y(n8236) );
  NAND2X1 U6675 ( .A(n8239), .B(n8240), .Y(n8238) );
  AOI21X1 U6676 ( .A0(n8240), .A1(n8241), .B0(test_se), .Y(n8237) );
  INVX1 U6677 ( .A(n8242), .Y(n8240) );
  AOI22X1 U6678 ( .A0(n8243), .A1(n8244), .B0(n13039), .B1(n7929), .Y(n8242)
         );
  AOI22X1 U6679 ( .A0(n8245), .A1(n13039), .B0(n13041), .B1(n7915), .Y(n8235)
         );
  NOR2X1 U6680 ( .A(n8246), .B(n7968), .Y(n8245) );
  OAI21X1 U6681 ( .A0(n7856), .A1(n7700), .B0(n8247), .Y(n7166) );
  AOI22X1 U6682 ( .A0(n8248), .A1(n8249), .B0(n12306), .B1(n8250), .Y(n8247)
         );
  OAI21X1 U6683 ( .A0(n7968), .A1(n8251), .B0(n8252), .Y(n8250) );
  AOI21X1 U6684 ( .A0(n8253), .A1(n8254), .B0(n8251), .Y(n8248) );
  MX2X1 U6685 ( .A(n8255), .B(n8256), .S0(n12303), .Y(n8254) );
  MX2X1 U6686 ( .A(n8257), .B(n8258), .S0(n7667), .Y(n8253) );
  OAI21X1 U6687 ( .A0(n7856), .A1(n7701), .B0(n8259), .Y(n7165) );
  AOI22X1 U6688 ( .A0(n8260), .A1(n8261), .B0(n12375), .B1(n8262), .Y(n8259)
         );
  OAI21X1 U6689 ( .A0(n7968), .A1(n8263), .B0(n8264), .Y(n8262) );
  AOI21X1 U6690 ( .A0(n8265), .A1(n8266), .B0(n8263), .Y(n8260) );
  MX2X1 U6691 ( .A(n8267), .B(n8268), .S0(n7660), .Y(n8266) );
  MX2X1 U6692 ( .A(n8269), .B(n8270), .S0(n12372), .Y(n8265) );
  OAI21X1 U6693 ( .A0(n12212), .A1(n8271), .B0(n8272), .Y(n7164) );
  AOI21X1 U6694 ( .A0(n8273), .A1(n12679), .B0(n8274), .Y(n8272) );
  AOI21X1 U6695 ( .A0(n7856), .A1(n8275), .B0(n7702), .Y(n8274) );
  NAND3X1 U6696 ( .A(n8276), .B(g35), .C(n12212), .Y(n8275) );
  NOR2X1 U6697 ( .A(n8276), .B(n7968), .Y(n8273) );
  AOI21X1 U6698 ( .A0(n8277), .A1(n8276), .B0(n7915), .Y(n8271) );
  NOR2X1 U6699 ( .A(test_se), .B(n12213), .Y(n8277) );
  OAI21X1 U6700 ( .A0(n7856), .A1(n7770), .B0(n8278), .Y(n7163) );
  AOI21X1 U6701 ( .A0(n12683), .A1(n7915), .B0(n8279), .Y(n8278) );
  AOI21X1 U6702 ( .A0(n8280), .A1(n7740), .B0(n7968), .Y(n8279) );
  OAI21X1 U6703 ( .A0(n12374), .A1(n7856), .B0(n8281), .Y(n7162) );
  AOI22X1 U6704 ( .A0(n8282), .A1(n3812), .B0(n12187), .B1(n7915), .Y(n8281)
         );
  NOR2X1 U6705 ( .A(n8283), .B(n7968), .Y(n8282) );
  AOI21X1 U6706 ( .A0(g9743), .A1(n7771), .B0(n12188), .Y(n8283) );
  OAI21X1 U6707 ( .A0(n12378), .A1(n7856), .B0(n8284), .Y(n7161) );
  AOI22X1 U6708 ( .A0(n8285), .A1(n3822), .B0(n12201), .B1(n7915), .Y(n8284)
         );
  NOR2X1 U6709 ( .A(n8286), .B(n7968), .Y(n8285) );
  AOI21X1 U6710 ( .A0(g9682), .A1(n7772), .B0(n12202), .Y(n8286) );
  OAI21X1 U6711 ( .A0(n12382), .A1(n7857), .B0(n8287), .Y(n7160) );
  AOI22X1 U6712 ( .A0(n8288), .A1(n3820), .B0(n12215), .B1(n7915), .Y(n8287)
         );
  NOR2X1 U6713 ( .A(n8289), .B(n7968), .Y(n8288) );
  AOI21X1 U6714 ( .A0(g9617), .A1(n7773), .B0(n12216), .Y(n8289) );
  OAI21X1 U6715 ( .A0(n12992), .A1(n7857), .B0(n8290), .Y(n7159) );
  AOI22X1 U6716 ( .A0(n8291), .A1(n3818), .B0(n12243), .B1(n7915), .Y(n8290)
         );
  NOR2X1 U6717 ( .A(n8292), .B(n7968), .Y(n8291) );
  AOI21X1 U6718 ( .A0(g9555), .A1(n7747), .B0(n12244), .Y(n8292) );
  OAI21X1 U6719 ( .A0(n12276), .A1(n7857), .B0(n8293), .Y(n7158) );
  AOI22X1 U6720 ( .A0(n8294), .A1(n3814), .B0(n12272), .B1(n7914), .Y(n8293)
         );
  NOR2X1 U6721 ( .A(n8295), .B(n7968), .Y(n8294) );
  AOI21X1 U6722 ( .A0(g9553), .A1(n7774), .B0(n12278), .Y(n8295) );
  OAI21X1 U6723 ( .A0(n7857), .A1(n7274), .B0(n8296), .Y(n7157) );
  AOI22X1 U6724 ( .A0(n8297), .A1(n3810), .B0(n12527), .B1(n7914), .Y(n8296)
         );
  NOR2X1 U6725 ( .A(n8298), .B(n7968), .Y(n8297) );
  AOI21X1 U6726 ( .A0(g8344), .A1(n7748), .B0(n12528), .Y(n8298) );
  OAI21X1 U6727 ( .A0(n7857), .A1(n7242), .B0(n8299), .Y(n7156) );
  AOI22X1 U6728 ( .A0(n8300), .A1(n7973), .B0(n12583), .B1(n7914), .Y(n8299)
         );
  NOR2X1 U6729 ( .A(n8301), .B(n7968), .Y(n8300) );
  AOI21X1 U6730 ( .A0(g8279), .A1(n7775), .B0(n12584), .Y(n8301) );
  OAI21X1 U6731 ( .A0(n7857), .A1(n7827), .B0(n8302), .Y(n7155) );
  AOI22X1 U6732 ( .A0(n8303), .A1(n7975), .B0(n12637), .B1(n7914), .Y(n8302)
         );
  NOR2X1 U6733 ( .A(n8304), .B(n7967), .Y(n8303) );
  AOI21X1 U6734 ( .A0(g8215), .A1(n7776), .B0(n12638), .Y(n8304) );
  OAI21X1 U6735 ( .A0(n7857), .A1(n7831), .B0(n8305), .Y(n7154) );
  AOI22X1 U6736 ( .A0(n12464), .A1(n7914), .B0(n12465), .B1(n7929), .Y(n8305)
         );
  OAI21X1 U6737 ( .A0(n8306), .A1(n7621), .B0(n8307), .Y(n7153) );
  NOR2X1 U6738 ( .A(n8308), .B(n8309), .Y(n8307) );
  AOI21X1 U6739 ( .A0(n7921), .A1(n8310), .B0(n12198), .Y(n8309) );
  NAND3X1 U6740 ( .A(n7668), .B(n7857), .C(n8311), .Y(n8310) );
  AOI21X1 U6741 ( .A0(n7857), .A1(n8312), .B0(n7668), .Y(n8308) );
  NAND3X1 U6742 ( .A(n8311), .B(g35), .C(n12198), .Y(n8312) );
  OAI21X1 U6743 ( .A0(n7857), .A1(n7287), .B0(n8313), .Y(n7152) );
  AOI22X1 U6744 ( .A0(n12754), .A1(n7914), .B0(n12750), .B1(n7929), .Y(n8313)
         );
  OAI21X1 U6745 ( .A0(n7857), .A1(n7466), .B0(n8314), .Y(n7151) );
  AOI22X1 U6746 ( .A0(n12763), .A1(n7914), .B0(n12751), .B1(n7929), .Y(n8314)
         );
  OAI21X1 U6747 ( .A0(n7857), .A1(n7290), .B0(n8315), .Y(n7150) );
  AOI22X1 U6748 ( .A0(n12781), .A1(n7914), .B0(n12778), .B1(n7929), .Y(n8315)
         );
  OAI21X1 U6749 ( .A0(n7857), .A1(n7294), .B0(n8316), .Y(n7149) );
  AOI22X1 U6750 ( .A0(n12833), .A1(n7914), .B0(n12830), .B1(n7929), .Y(n8316)
         );
  OAI21X1 U6751 ( .A0(n7857), .A1(n7292), .B0(n8317), .Y(n7148) );
  AOI22X1 U6752 ( .A0(n12857), .A1(n7914), .B0(n12854), .B1(n7929), .Y(n8317)
         );
  OAI21X1 U6753 ( .A0(n7858), .A1(n7470), .B0(n8318), .Y(n7147) );
  AOI22X1 U6754 ( .A0(n12867), .A1(n7914), .B0(n12855), .B1(n7929), .Y(n8318)
         );
  OAI21X1 U6755 ( .A0(n7858), .A1(n7404), .B0(n8319), .Y(n7146) );
  AOI22X1 U6756 ( .A0(n12879), .A1(n7914), .B0(n12876), .B1(n7929), .Y(n8319)
         );
  OAI21X1 U6757 ( .A0(n7858), .A1(n7421), .B0(n8320), .Y(n7145) );
  AOI22X1 U6758 ( .A0(n12889), .A1(n7913), .B0(n12877), .B1(n7929), .Y(n8320)
         );
  OAI21X1 U6759 ( .A0(n7858), .A1(n7777), .B0(n8321), .Y(n7144) );
  AOI22X1 U6760 ( .A0(n12469), .A1(n7913), .B0(n12464), .B1(n7929), .Y(n8321)
         );
  OAI21X1 U6761 ( .A0(n7858), .A1(n7339), .B0(n8322), .Y(n7143) );
  AOI22X1 U6762 ( .A0(n12473), .A1(n7913), .B0(n12471), .B1(n7929), .Y(n8322)
         );
  OAI21X1 U6763 ( .A0(n7858), .A1(n7759), .B0(n8323), .Y(n7142) );
  AOI22X1 U6764 ( .A0(n12639), .A1(n7913), .B0(n12640), .B1(n7929), .Y(n8323)
         );
  OAI21X1 U6765 ( .A0(n7858), .A1(n7832), .B0(n8324), .Y(n7141) );
  AOI22X1 U6766 ( .A0(n12680), .A1(n7913), .B0(n12661), .B1(n7929), .Y(n8324)
         );
  OAI21X1 U6767 ( .A0(n7858), .A1(n7740), .B0(n8325), .Y(n7140) );
  AOI22X1 U6768 ( .A0(n12682), .A1(n7913), .B0(n12680), .B1(n7929), .Y(n8325)
         );
  OAI21X1 U6769 ( .A0(n7858), .A1(n7741), .B0(n8326), .Y(n7139) );
  AOI22X1 U6770 ( .A0(n12685), .A1(n7913), .B0(n12682), .B1(n7929), .Y(n8326)
         );
  OAI21X1 U6771 ( .A0(n7858), .A1(g23652), .B0(n8327), .Y(n7138) );
  AOI22X1 U6772 ( .A0(n12684), .A1(n7913), .B0(n12685), .B1(n7929), .Y(n8327)
         );
  OAI21X1 U6773 ( .A0(n7858), .A1(n7468), .B0(n8328), .Y(n7137) );
  AOI22X1 U6774 ( .A0(n12721), .A1(n7913), .B0(n12709), .B1(n7929), .Y(n8328)
         );
  OAI21X1 U6775 ( .A0(n7858), .A1(n7467), .B0(n8329), .Y(n7136) );
  AOI22X1 U6776 ( .A0(n12742), .A1(n7913), .B0(n12730), .B1(n7929), .Y(n8329)
         );
  OAI21X1 U6777 ( .A0(n7858), .A1(n7465), .B0(n8330), .Y(n7135) );
  AOI22X1 U6778 ( .A0(n12792), .A1(n7913), .B0(n12779), .B1(n7929), .Y(n8330)
         );
  OAI21X1 U6779 ( .A0(n7858), .A1(n7293), .B0(n8331), .Y(n7134) );
  AOI22X1 U6780 ( .A0(n12843), .A1(n7913), .B0(n12831), .B1(n7929), .Y(n8331)
         );
  OAI21X1 U6781 ( .A0(n7858), .A1(n7778), .B0(n8332), .Y(n7133) );
  AOI22X1 U6782 ( .A0(n8333), .A1(n12523), .B0(n12300), .B1(n8334), .Y(n8332)
         );
  OAI21X1 U6783 ( .A0(test_se), .A1(n8335), .B0(n7918), .Y(n8334) );
  AND2X1 U6784 ( .A(n8335), .B(n7929), .Y(n8333) );
  OAI21X1 U6785 ( .A0(n7858), .A1(n7285), .B0(n8336), .Y(n7132) );
  AOI22X1 U6786 ( .A0(n8337), .A1(n12391), .B0(n12306), .B1(n8338), .Y(n8336)
         );
  OAI21X1 U6787 ( .A0(test_se), .A1(n8251), .B0(n7918), .Y(n8338) );
  AND2X1 U6788 ( .A(n8251), .B(n7929), .Y(n8337) );
  NAND2X1 U6789 ( .A(n8339), .B(n8340), .Y(n8251) );
  OAI21X1 U6790 ( .A0(n7858), .A1(n7669), .B0(n8341), .Y(n7131) );
  AOI22X1 U6791 ( .A0(n8342), .A1(n12400), .B0(n12375), .B1(n8343), .Y(n8341)
         );
  OAI21X1 U6792 ( .A0(test_se), .A1(n8263), .B0(n7918), .Y(n8343) );
  AND2X1 U6793 ( .A(n8263), .B(n7929), .Y(n8342) );
  NAND2X1 U6794 ( .A(n8344), .B(n8345), .Y(n8263) );
  NAND2X1 U6795 ( .A(n8346), .B(n8347), .Y(n7130) );
  AOI22X1 U6796 ( .A0(n8249), .A1(n8348), .B0(n12299), .B1(n7910), .Y(n8347)
         );
  AOI22X1 U6797 ( .A0(n8349), .A1(n12387), .B0(test_se), .B1(n7411), .Y(n8346)
         );
  NAND2X1 U6798 ( .A(n8350), .B(n8351), .Y(n7129) );
  AOI22X1 U6799 ( .A0(n8352), .A1(n8353), .B0(n8215), .B1(n12396), .Y(n8351)
         );
  AOI22X1 U6800 ( .A0(n12327), .A1(n7910), .B0(test_se), .B1(n7504), .Y(n8350)
         );
  NAND2X1 U6801 ( .A(n8354), .B(n8355), .Y(n7128) );
  AOI22X1 U6802 ( .A0(n8356), .A1(n8357), .B0(n12394), .B1(n8358), .Y(n8355)
         );
  AND2X1 U6803 ( .A(n7930), .B(n8359), .Y(n8356) );
  AOI22X1 U6804 ( .A0(n12371), .A1(n7910), .B0(test_se), .B1(n7255), .Y(n8354)
         );
  NAND2X1 U6805 ( .A(n8360), .B(n8361), .Y(n7127) );
  AOI22X1 U6806 ( .A0(n8362), .A1(n8199), .B0(n8363), .B1(n12531), .Y(n8361)
         );
  AOI22X1 U6807 ( .A0(n12554), .A1(n7910), .B0(n12566), .B1(test_se), .Y(n8360) );
  NAND2X1 U6808 ( .A(n8364), .B(n8365), .Y(n7126) );
  AOI22X1 U6809 ( .A0(n8366), .A1(n7930), .B0(n8367), .B1(n12707), .Y(n8365)
         );
  AOI21X1 U6810 ( .A0(n8368), .A1(n8369), .B0(n8370), .Y(n8366) );
  AOI21X1 U6811 ( .A0(n12707), .A1(n8371), .B0(n8372), .Y(n8370) );
  INVX1 U6812 ( .A(n8373), .Y(n8369) );
  INVX1 U6813 ( .A(n8374), .Y(n8368) );
  AOI21X1 U6814 ( .A0(n8372), .A1(n12707), .B0(n8375), .Y(n8374) );
  OR2X1 U6815 ( .A(n7529), .B(n8376), .Y(n8372) );
  AOI22X1 U6816 ( .A0(n12722), .A1(n7910), .B0(n13023), .B1(test_se), .Y(n8364) );
  NAND2X1 U6817 ( .A(n8377), .B(n8378), .Y(n7125) );
  AOI22X1 U6818 ( .A0(n8379), .A1(n7930), .B0(n8380), .B1(n12728), .Y(n8378)
         );
  AOI21X1 U6819 ( .A0(n8381), .A1(n8382), .B0(n8383), .Y(n8379) );
  AOI21X1 U6820 ( .A0(n12728), .A1(n8384), .B0(n8385), .Y(n8383) );
  INVX1 U6821 ( .A(n8386), .Y(n8382) );
  INVX1 U6822 ( .A(n8387), .Y(n8381) );
  AOI21X1 U6823 ( .A0(n8385), .A1(n12728), .B0(n8388), .Y(n8387) );
  NAND2X1 U6824 ( .A(n8389), .B(n7529), .Y(n8385) );
  AOI22X1 U6825 ( .A0(n12743), .A1(n7910), .B0(n13024), .B1(test_se), .Y(n8377) );
  NAND2X1 U6826 ( .A(n8390), .B(n8391), .Y(n7124) );
  AOI22X1 U6827 ( .A0(n8392), .A1(n7930), .B0(n8393), .B1(n12749), .Y(n8391)
         );
  AOI21X1 U6828 ( .A0(n8394), .A1(n8395), .B0(n8396), .Y(n8392) );
  AOI21X1 U6829 ( .A0(n12749), .A1(n8397), .B0(n8398), .Y(n8396) );
  INVX1 U6830 ( .A(n8399), .Y(n8395) );
  INVX1 U6831 ( .A(n8400), .Y(n8394) );
  AOI21X1 U6832 ( .A0(n8398), .A1(n12749), .B0(n8401), .Y(n8400) );
  NAND2X1 U6833 ( .A(n8402), .B(n12895), .Y(n8398) );
  AOI22X1 U6834 ( .A0(n12764), .A1(n7910), .B0(n13022), .B1(test_se), .Y(n8390) );
  NAND2X1 U6835 ( .A(n8403), .B(n8404), .Y(n7123) );
  AOI21X1 U6836 ( .A0(n8405), .A1(n12776), .B0(n8406), .Y(n8404) );
  AOI21X1 U6837 ( .A0(n8407), .A1(n8408), .B0(n8409), .Y(n8406) );
  AOI21X1 U6838 ( .A0(n8410), .A1(n7930), .B0(n8411), .Y(n8409) );
  AOI21X1 U6839 ( .A0(n12776), .A1(n8412), .B0(n8413), .Y(n8410) );
  INVX1 U6840 ( .A(n8407), .Y(n8412) );
  OAI21X1 U6841 ( .A0(n12793), .A1(n12792), .B0(n12776), .Y(n8408) );
  NOR2X1 U6842 ( .A(n8414), .B(n12895), .Y(n8407) );
  AOI22X1 U6843 ( .A0(n12793), .A1(n7910), .B0(n13025), .B1(test_se), .Y(n8403) );
  OAI21X1 U6844 ( .A0(n7858), .A1(n7315), .B0(n8415), .Y(n7122) );
  AOI22X1 U6845 ( .A0(n7930), .A1(n8416), .B0(n12820), .B1(n7910), .Y(n8415)
         );
  INVX1 U6846 ( .A(n8417), .Y(n8416) );
  AOI22X1 U6847 ( .A0(n8418), .A1(n8419), .B0(n8420), .B1(n12799), .Y(n8417)
         );
  INVX1 U6848 ( .A(n8421), .Y(n8420) );
  AOI21X1 U6849 ( .A0(n8422), .A1(n8418), .B0(n8423), .Y(n8421) );
  OR2X1 U6850 ( .A(n8424), .B(n8425), .Y(n8418) );
  AOI21X1 U6851 ( .A0(n12799), .A1(n8419), .B0(n8423), .Y(n8425) );
  NAND2X1 U6852 ( .A(n8426), .B(n13035), .Y(n8419) );
  NAND2X1 U6853 ( .A(n8427), .B(n8428), .Y(n7121) );
  AOI22X1 U6854 ( .A0(n8429), .A1(n8430), .B0(n8431), .B1(n12826), .Y(n8428)
         );
  OAI21X1 U6855 ( .A0(n8432), .A1(n8433), .B0(n8434), .Y(n8430) );
  INVX1 U6856 ( .A(n8435), .Y(n8434) );
  AOI21X1 U6857 ( .A0(n8436), .A1(n7282), .B0(n7703), .Y(n8432) );
  OAI21X1 U6858 ( .A0(n8437), .A1(n7967), .B0(n8438), .Y(n8429) );
  AOI21X1 U6859 ( .A0(n12826), .A1(n8439), .B0(n8440), .Y(n8437) );
  AOI22X1 U6860 ( .A0(n12844), .A1(n7910), .B0(n13014), .B1(test_se), .Y(n8427) );
  OAI21X1 U6861 ( .A0(n7858), .A1(n7524), .B0(n8441), .Y(n7120) );
  AOI22X1 U6862 ( .A0(n7930), .A1(n8442), .B0(n12868), .B1(n7910), .Y(n8441)
         );
  INVX1 U6863 ( .A(n8443), .Y(n8442) );
  AOI22X1 U6864 ( .A0(n8444), .A1(n8445), .B0(n8446), .B1(n12853), .Y(n8443)
         );
  INVX1 U6865 ( .A(n8447), .Y(n8446) );
  AOI21X1 U6866 ( .A0(n8448), .A1(n8444), .B0(n8449), .Y(n8447) );
  OR2X1 U6867 ( .A(n8450), .B(n8451), .Y(n8444) );
  AOI21X1 U6868 ( .A0(n12853), .A1(n8445), .B0(n8449), .Y(n8451) );
  NAND2X1 U6869 ( .A(n8426), .B(n7367), .Y(n8445) );
  AND2X1 U6870 ( .A(n8452), .B(n7500), .Y(n8426) );
  NAND2X1 U6871 ( .A(n8453), .B(n8454), .Y(n7119) );
  AOI22X1 U6872 ( .A0(n8455), .A1(n7930), .B0(n8456), .B1(n12875), .Y(n8454)
         );
  AOI21X1 U6873 ( .A0(n8457), .A1(n8436), .B0(n8458), .Y(n8455) );
  AOI21X1 U6874 ( .A0(n8459), .A1(n8460), .B0(n8461), .Y(n8458) );
  OAI21X1 U6875 ( .A0(n13041), .A1(n8440), .B0(n12875), .Y(n8459) );
  INVX1 U6876 ( .A(n8440), .Y(n8436) );
  NAND2X1 U6877 ( .A(n13006), .B(n8452), .Y(n8440) );
  AOI21X1 U6878 ( .A0(n12875), .A1(n8462), .B0(n13041), .Y(n8457) );
  AOI22X1 U6879 ( .A0(n12890), .A1(n7910), .B0(n13015), .B1(test_se), .Y(n8453) );
  NAND2X1 U6880 ( .A(n8463), .B(n8464), .Y(n7118) );
  AOI22X1 U6881 ( .A0(n8465), .A1(n8466), .B0(n8467), .B1(n12970), .Y(n8464)
         );
  AOI21X1 U6882 ( .A0(n8468), .A1(n8466), .B0(n7967), .Y(n8467) );
  NOR2X1 U6883 ( .A(n8468), .B(n8469), .Y(n8465) );
  XOR2X1 U6884 ( .A(n8230), .B(n7534), .Y(n8468) );
  AOI22X1 U6885 ( .A0(n12908), .A1(n7909), .B0(n12913), .B1(test_se), .Y(n8463) );
  NAND2X1 U6886 ( .A(n8470), .B(n8471), .Y(n7117) );
  AOI22X1 U6887 ( .A0(n8472), .A1(n8473), .B0(n13034), .B1(n8474), .Y(n8471)
         );
  XOR2X1 U6888 ( .A(n8239), .B(n7362), .Y(n8473) );
  AOI21X1 U6889 ( .A0(n7611), .A1(n8475), .B0(n7967), .Y(n8472) );
  NAND3X1 U6890 ( .A(n7272), .B(n7679), .C(n8476), .Y(n8475) );
  AOI22X1 U6891 ( .A0(n13036), .A1(n7909), .B0(n13041), .B1(test_se), .Y(n8470) );
  NAND2X1 U6892 ( .A(n8477), .B(n8478), .Y(n7116) );
  AOI22X1 U6893 ( .A0(n8479), .A1(n8480), .B0(n12328), .B1(n8481), .Y(n8478)
         );
  AOI22X1 U6894 ( .A0(n12920), .A1(n7909), .B0(n12178), .B1(test_se), .Y(n8477) );
  OAI21X1 U6895 ( .A0(n12198), .A1(n7858), .B0(n8482), .Y(n7115) );
  AOI22X1 U6896 ( .A0(n12195), .A1(n8483), .B0(n8484), .B1(n12199), .Y(n8482)
         );
  OAI21X1 U6897 ( .A0(test_se), .A1(n8485), .B0(n7918), .Y(n8483) );
  OAI21X1 U6898 ( .A0(n12212), .A1(n7858), .B0(n8486), .Y(n7114) );
  AOI22X1 U6899 ( .A0(n12209), .A1(n8487), .B0(n8488), .B1(n12213), .Y(n8486)
         );
  OAI21X1 U6900 ( .A0(test_se), .A1(n8489), .B0(n7918), .Y(n8487) );
  OAI21X1 U6901 ( .A0(n12239), .A1(n7858), .B0(n8490), .Y(n7113) );
  AOI22X1 U6902 ( .A0(n12235), .A1(n8491), .B0(n12238), .B1(n8492), .Y(n8490)
         );
  OAI21X1 U6903 ( .A0(test_se), .A1(n8493), .B0(n7918), .Y(n8491) );
  OAI21X1 U6904 ( .A0(n12257), .A1(n7858), .B0(n8494), .Y(n7112) );
  AOI22X1 U6905 ( .A0(n12254), .A1(n8495), .B0(n12258), .B1(n8496), .Y(n8494)
         );
  OAI21X1 U6906 ( .A0(test_se), .A1(n8497), .B0(n7918), .Y(n8495) );
  OAI21X1 U6907 ( .A0(n7858), .A1(n7513), .B0(n8498), .Y(n7111) );
  AOI22X1 U6908 ( .A0(n12497), .A1(n8499), .B0(n12500), .B1(n8500), .Y(n8498)
         );
  OAI21X1 U6909 ( .A0(test_se), .A1(n8501), .B0(n7918), .Y(n8499) );
  OAI21X1 U6910 ( .A0(n7859), .A1(n7526), .B0(n8502), .Y(n7110) );
  AOI22X1 U6911 ( .A0(n12545), .A1(n8503), .B0(n12548), .B1(n8504), .Y(n8502)
         );
  OAI21X1 U6912 ( .A0(test_se), .A1(n8505), .B0(n7918), .Y(n8503) );
  OAI21X1 U6913 ( .A0(n12602), .A1(n7859), .B0(n8506), .Y(n7109) );
  AOI22X1 U6914 ( .A0(n12599), .A1(n8507), .B0(n12634), .B1(n8508), .Y(n8506)
         );
  INVX1 U6915 ( .A(n8509), .Y(n8507) );
  AOI21X1 U6916 ( .A0(n7859), .A1(n8510), .B0(n7909), .Y(n8509) );
  NAND2X1 U6917 ( .A(n8511), .B(n8512), .Y(n7108) );
  AOI22X1 U6918 ( .A0(n12457), .A1(n8513), .B0(n8514), .B1(n7205), .Y(n8512)
         );
  AOI22X1 U6919 ( .A0(n12476), .A1(n7909), .B0(n12487), .B1(test_se), .Y(n8511) );
  OAI21X1 U6920 ( .A0(n7859), .A1(n7704), .B0(n8515), .Y(n7107) );
  AOI22X1 U6921 ( .A0(n8516), .A1(n8517), .B0(n12300), .B1(n8518), .Y(n8515)
         );
  OAI21X1 U6922 ( .A0(n7967), .A1(n8335), .B0(n8519), .Y(n8518) );
  INVX1 U6923 ( .A(n8520), .Y(n8519) );
  AOI21X1 U6924 ( .A0(n8521), .A1(n8522), .B0(n8335), .Y(n8516) );
  NAND2X1 U6925 ( .A(n8339), .B(n8523), .Y(n8335) );
  MX2X1 U6926 ( .A(n8524), .B(n8525), .S0(n12485), .Y(n8522) );
  MX2X1 U6927 ( .A(n8526), .B(n8527), .S0(n12484), .Y(n8521) );
  INVX1 U6928 ( .A(n8528), .Y(n7106) );
  AOI21X1 U6929 ( .A0(n8529), .A1(n8530), .B0(n8531), .Y(n8528) );
  MX2X1 U6930 ( .A(n12267), .B(n12926), .S0(n8532), .Y(n8531) );
  OAI21X1 U6931 ( .A0(n7859), .A1(n7642), .B0(n8533), .Y(n7105) );
  MX2X1 U6932 ( .A(n8534), .B(n8535), .S0(n8536), .Y(n8533) );
  AND2X1 U6933 ( .A(n8485), .B(n12195), .Y(n8536) );
  INVX1 U6934 ( .A(n8537), .Y(n8485) );
  OAI21X1 U6935 ( .A0(n7859), .A1(n7641), .B0(n8538), .Y(n7104) );
  MX2X1 U6936 ( .A(n8534), .B(n8535), .S0(n8539), .Y(n8538) );
  AND2X1 U6937 ( .A(n8489), .B(n12209), .Y(n8539) );
  INVX1 U6938 ( .A(n8540), .Y(n8489) );
  OAI21X1 U6939 ( .A0(n7854), .A1(n7622), .B0(n8541), .Y(n7103) );
  MX2X1 U6940 ( .A(n8534), .B(n8535), .S0(n8542), .Y(n8541) );
  AND2X1 U6941 ( .A(n8493), .B(n12235), .Y(n8542) );
  INVX1 U6942 ( .A(n8543), .Y(n8493) );
  OAI21X1 U6943 ( .A0(n7859), .A1(n7646), .B0(n8544), .Y(n7102) );
  MX2X1 U6944 ( .A(n8534), .B(n8535), .S0(n8545), .Y(n8544) );
  AND2X1 U6945 ( .A(n8497), .B(n12254), .Y(n8545) );
  INVX1 U6946 ( .A(g32975), .Y(n8497) );
  OAI21X1 U6947 ( .A0(n7859), .A1(n7334), .B0(n8546), .Y(n7101) );
  MX2X1 U6948 ( .A(n8534), .B(n8535), .S0(n8547), .Y(n8546) );
  AND2X1 U6949 ( .A(n8501), .B(n12497), .Y(n8547) );
  INVX1 U6950 ( .A(n8548), .Y(n8501) );
  OAI21X1 U6951 ( .A0(n7859), .A1(n7333), .B0(n8549), .Y(n7100) );
  MX2X1 U6952 ( .A(n8534), .B(n8535), .S0(n8550), .Y(n8549) );
  AND2X1 U6953 ( .A(n8505), .B(n12545), .Y(n8550) );
  INVX1 U6954 ( .A(n8551), .Y(n8505) );
  OAI21X1 U6955 ( .A0(n7859), .A1(n7644), .B0(n8552), .Y(n7099) );
  MX2X1 U6956 ( .A(n8534), .B(n8535), .S0(n8553), .Y(n8552) );
  NOR2X1 U6957 ( .A(n8510), .B(n7745), .Y(n8553) );
  OAI21X1 U6958 ( .A0(n7859), .A1(n7323), .B0(n8554), .Y(n7098) );
  MX2X1 U6959 ( .A(n8534), .B(n8535), .S0(n8555), .Y(n8554) );
  AND2X1 U6960 ( .A(n8556), .B(n12180), .Y(n8555) );
  NAND2X1 U6961 ( .A(n8557), .B(n7930), .Y(n8535) );
  OAI21X1 U6962 ( .A0(n7859), .A1(n7321), .B0(n8558), .Y(n7097) );
  AOI22X1 U6963 ( .A0(n12457), .A1(n8559), .B0(n12487), .B1(n8513), .Y(n8558)
         );
  OAI21X1 U6964 ( .A0(n7859), .A1(n7756), .B0(n8560), .Y(n7096) );
  AOI22X1 U6965 ( .A0(n12925), .A1(n8561), .B0(n8562), .B1(n12924), .Y(n8560)
         );
  OAI21X1 U6966 ( .A0(test_se), .A1(n8563), .B0(n7918), .Y(n8561) );
  INVX1 U6967 ( .A(n8564), .Y(n7094) );
  MX2X1 U6968 ( .A(n7975), .B(n489), .S0(n8104), .Y(n8564) );
  MX2X1 U6969 ( .A(g16718), .B(g14421), .S0(n8104), .Y(n7093) );
  INVX1 U6970 ( .A(n8565), .Y(n7092) );
  MX2X1 U6971 ( .A(n7973), .B(n524), .S0(n8104), .Y(n8565) );
  MX2X1 U6972 ( .A(g16744), .B(g14451), .S0(n8104), .Y(n7091) );
  INVX1 U6973 ( .A(n8566), .Y(n7090) );
  MX2X1 U6974 ( .A(n3810), .B(n7984), .S0(n8104), .Y(n8566) );
  MX2X1 U6975 ( .A(g16775), .B(g14518), .S0(n8104), .Y(n7089) );
  INVX1 U6976 ( .A(n8567), .Y(n7088) );
  MX2X1 U6977 ( .A(n7826), .B(n5243), .S0(n8104), .Y(n8567) );
  INVX1 U6978 ( .A(n8568), .Y(n7087) );
  MX2X1 U6979 ( .A(n5243), .B(n5242), .S0(n8104), .Y(n8568) );
  MX2X1 U6980 ( .A(n12429), .B(n12426), .S0(n7865), .Y(n7086) );
  MX2X1 U6981 ( .A(n12449), .B(n12427), .S0(n7868), .Y(n7085) );
  MX2X1 U6982 ( .A(n12423), .B(n12416), .S0(n7854), .Y(n7084) );
  MX2X1 U6983 ( .A(n12407), .B(n12157), .S0(n7846), .Y(n7083) );
  MX2X1 U6984 ( .A(g9553), .B(g9497), .S0(n7845), .Y(n7082) );
  MX2X1 U6985 ( .A(n12266), .B(g9553), .S0(n7847), .Y(n7081) );
  MX2X1 U6986 ( .A(g17674), .B(g13039), .S0(n7849), .Y(n7080) );
  INVX1 U6987 ( .A(n8569), .Y(n7079) );
  MX2X1 U6988 ( .A(n3818), .B(n7990), .S0(n7848), .Y(n8569) );
  MX2X1 U6989 ( .A(g17711), .B(g13049), .S0(n7851), .Y(n7078) );
  INVX1 U6990 ( .A(n8570), .Y(n7077) );
  MX2X1 U6991 ( .A(n3820), .B(n7992), .S0(n7852), .Y(n8570) );
  MX2X1 U6992 ( .A(g17739), .B(g13068), .S0(n7853), .Y(n7076) );
  INVX1 U6993 ( .A(n8571), .Y(n7075) );
  MX2X1 U6994 ( .A(n3822), .B(n7994), .S0(n7845), .Y(n8571) );
  MX2X1 U6995 ( .A(g17760), .B(g13085), .S0(n7845), .Y(n7074) );
  INVX1 U6996 ( .A(n8572), .Y(n7073) );
  MX2X1 U6997 ( .A(n3812), .B(n7986), .S0(n7845), .Y(n8572) );
  MX2X1 U6998 ( .A(g17778), .B(g13099), .S0(n7845), .Y(n7072) );
  MX2X1 U6999 ( .A(n12159), .B(g11678), .S0(n7845), .Y(n7071) );
  MX2X1 U7000 ( .A(n12769), .B(g14189), .S0(n7845), .Y(n7070) );
  MX2X1 U7001 ( .A(g14201), .B(g14167), .S0(n7845), .Y(n7069) );
  MX2X1 U7002 ( .A(n12772), .B(g14201), .S0(n7846), .Y(n7068) );
  INVX1 U7003 ( .A(n8573), .Y(n7067) );
  AOI22X1 U7004 ( .A0(n7909), .A1(n7385), .B0(n12228), .B1(test_se), .Y(n8573)
         );
  INVX1 U7005 ( .A(n8574), .Y(n7066) );
  AOI22X1 U7006 ( .A0(n12814), .A1(n7909), .B0(n12812), .B1(test_se), .Y(n8574) );
  MX2X1 U7007 ( .A(n12386), .B(g4549), .S0(n8155), .Y(n7065) );
  MX2X1 U7008 ( .A(n12393), .B(g4504), .S0(n8155), .Y(n7064) );
  INVX1 U7009 ( .A(n8575), .Y(n7063) );
  AOI22X1 U7010 ( .A0(n7930), .A1(g21176), .B0(n12489), .B1(test_se), .Y(n8575) );
  OAI21X1 U7011 ( .A0(n7857), .A1(n7779), .B0(n8576), .Y(n7062) );
  AOI22X1 U7012 ( .A0(n8577), .A1(n12550), .B0(n12301), .B1(n8578), .Y(n8576)
         );
  OAI21X1 U7013 ( .A0(test_se), .A1(n8201), .B0(n7918), .Y(n8578) );
  AND2X1 U7014 ( .A(n8201), .B(n7930), .Y(n8577) );
  NAND2X1 U7015 ( .A(n8339), .B(n8579), .Y(n8201) );
  OAI21X1 U7016 ( .A0(n7857), .A1(n7780), .B0(n8580), .Y(n7061) );
  AOI22X1 U7017 ( .A0(n8581), .A1(n12402), .B0(n12379), .B1(n8582), .Y(n8580)
         );
  INVX1 U7018 ( .A(n8583), .Y(n8582) );
  AOI21X1 U7019 ( .A0(n7857), .A1(n8214), .B0(n7909), .Y(n8583) );
  NOR2X1 U7020 ( .A(n8214), .B(n7967), .Y(n8581) );
  NOR2X1 U7021 ( .A(n8584), .B(n8585), .Y(n8214) );
  INVX1 U7022 ( .A(n8586), .Y(n7060) );
  AOI22X1 U7023 ( .A0(n7930), .A1(n8587), .B0(test_se), .B1(n7353), .Y(n8586)
         );
  NAND4X1 U7024 ( .A(n8139), .B(n8588), .C(n8589), .D(n7412), .Y(n8587) );
  NOR2X1 U7025 ( .A(n12451), .B(n12452), .Y(n8589) );
  INVX1 U7026 ( .A(n8590), .Y(n7059) );
  AOI22X1 U7027 ( .A0(n7930), .A1(n7623), .B0(n12462), .B1(test_se), .Y(n8590)
         );
  MX2X1 U7028 ( .A(n8591), .B(n8592), .S0(n7650), .Y(n7058) );
  NOR2X1 U7029 ( .A(n5244), .B(n7967), .Y(n8592) );
  OR2X1 U7030 ( .A(n8593), .B(n5244), .Y(n8591) );
  INVX1 U7031 ( .A(n8594), .Y(n7057) );
  AOI22X1 U7032 ( .A0(n7930), .A1(n7625), .B0(n12469), .B1(test_se), .Y(n8594)
         );
  MX2X1 U7033 ( .A(g18095), .B(n12412), .S0(n7959), .Y(n7056) );
  MX2X1 U7034 ( .A(g18094), .B(n12413), .S0(n7959), .Y(n7055) );
  MX2X1 U7035 ( .A(g18096), .B(n12421), .S0(n7958), .Y(n7054) );
  MX2X1 U7036 ( .A(g18095), .B(n12420), .S0(n7958), .Y(n7053) );
  MX2X1 U7037 ( .A(g18094), .B(n12419), .S0(n7958), .Y(n7052) );
  MX2X1 U7038 ( .A(n7539), .B(n12593), .S0(n7958), .Y(n7051) );
  MX2X1 U7039 ( .A(n8595), .B(n7967), .S0(n12158), .Y(n7050) );
  AOI21X1 U7040 ( .A0(n7705), .A1(n7342), .B0(n7967), .Y(n8595) );
  MX2X1 U7041 ( .A(n8596), .B(n12641), .S0(n7957), .Y(n7049) );
  NAND2X1 U7042 ( .A(n12536), .B(n7743), .Y(n8596) );
  MX2X1 U7043 ( .A(n12829), .B(n12892), .S0(n7957), .Y(n7048) );
  MX2X1 U7044 ( .A(n12157), .B(n8185), .S0(n7846), .Y(n7046) );
  AND2X1 U7045 ( .A(g35), .B(n8597), .Y(n8185) );
  NAND2X1 U7046 ( .A(n8598), .B(n8599), .Y(n8597) );
  AOI22X1 U7047 ( .A0(n4770), .A1(n7781), .B0(n12531), .B1(n4771), .Y(n8599)
         );
  AOI21X1 U7048 ( .A0(n12387), .A1(n7431), .B0(n8600), .Y(n8598) );
  MX2X1 U7049 ( .A(n7782), .B(n8601), .S0(n7285), .Y(n8600) );
  AOI21X1 U7050 ( .A0(n8602), .A1(n8603), .B0(n8604), .Y(n8601) );
  MX2X1 U7051 ( .A(n8605), .B(n8606), .S0(n7250), .Y(n8602) );
  NAND2X1 U7052 ( .A(n12610), .B(n8607), .Y(n8606) );
  NAND2X1 U7053 ( .A(n12608), .B(n8608), .Y(n8605) );
  MX2X1 U7054 ( .A(n8609), .B(n8610), .S0(n7363), .Y(n8608) );
  INVX1 U7055 ( .A(n8611), .Y(n8610) );
  XOR2X1 U7056 ( .A(n8612), .B(n8607), .Y(n8611) );
  NAND2X1 U7057 ( .A(n8613), .B(n8614), .Y(n8607) );
  AOI22X1 U7058 ( .A0(n8579), .A1(n7499), .B0(n12523), .B1(n8340), .Y(n8614)
         );
  AOI22X1 U7059 ( .A0(n12550), .A1(n8523), .B0(n12391), .B1(n8615), .Y(n8613)
         );
  AOI22X1 U7060 ( .A0(n12390), .A1(n8579), .B0(n12389), .B1(n8615), .Y(n8612)
         );
  NAND3X1 U7061 ( .A(n8616), .B(n8617), .C(n8618), .Y(n8609) );
  NAND2X1 U7062 ( .A(n8340), .B(n7746), .Y(n8618) );
  INVX1 U7063 ( .A(n8523), .Y(n8617) );
  MX2X1 U7064 ( .A(n12536), .B(n8188), .S0(n7846), .Y(n7045) );
  AND2X1 U7065 ( .A(g35), .B(n8619), .Y(n8188) );
  NAND2X1 U7066 ( .A(n8620), .B(n8621), .Y(n8619) );
  AOI22X1 U7067 ( .A0(n12995), .A1(g21245), .B0(n6763), .B1(n7783), .Y(n8621)
         );
  AOI21X1 U7068 ( .A0(n12396), .A1(n4749), .B0(n8622), .Y(n8620) );
  MX2X1 U7069 ( .A(n8623), .B(n12395), .S0(n7360), .Y(n8622) );
  AOI21X1 U7070 ( .A0(n8584), .A1(n8624), .B0(n8625), .Y(n8623) );
  NAND2X1 U7071 ( .A(n8626), .B(n8627), .Y(n8624) );
  OAI21X1 U7072 ( .A0(n8628), .A1(n7354), .B0(n7246), .Y(n8627) );
  XOR2X1 U7073 ( .A(n8629), .B(n8630), .Y(n8628) );
  AOI22X1 U7074 ( .A0(n12398), .A1(n8631), .B0(n12397), .B1(n8632), .Y(n8630)
         );
  MX2X1 U7075 ( .A(n8633), .B(n8629), .S0(n7354), .Y(n8626) );
  NAND2X1 U7076 ( .A(n8634), .B(n8635), .Y(n8629) );
  AOI22X1 U7077 ( .A0(n8631), .A1(n7442), .B0(n12402), .B1(n8345), .Y(n8635)
         );
  AOI22X1 U7078 ( .A0(n12400), .A1(n8636), .B0(n13002), .B1(n8632), .Y(n8634)
         );
  AOI21X1 U7079 ( .A0(n8637), .A1(n8638), .B0(n7255), .Y(n8633) );
  NOR2X1 U7080 ( .A(n8345), .B(n8631), .Y(n8638) );
  AOI21X1 U7081 ( .A0(n8636), .A1(n7751), .B0(n7246), .Y(n8637) );
  NAND2X1 U7082 ( .A(n8639), .B(n8640), .Y(n6865) );
  MX2X1 U7083 ( .A(n671), .B(n8641), .S0(n7846), .Y(n8640) );
  NAND2X1 U7084 ( .A(n8642), .B(n7573), .Y(n8641) );
  AOI22X1 U7085 ( .A0(n12228), .A1(n7909), .B0(n8643), .B1(n8562), .Y(n8639)
         );
  NOR2X1 U7086 ( .A(n8642), .B(n7573), .Y(n8643) );
  INVX1 U7087 ( .A(n8563), .Y(n8642) );
  NAND2X1 U7088 ( .A(n12228), .B(n8644), .Y(n8563) );
  NAND2X1 U7089 ( .A(n8645), .B(n8646), .Y(n6864) );
  MX2X1 U7090 ( .A(n7316), .B(n8647), .S0(n7846), .Y(n8646) );
  NAND3X1 U7091 ( .A(n8648), .B(n7607), .C(n8649), .Y(n8647) );
  AOI22X1 U7092 ( .A0(n12904), .A1(n7909), .B0(n8650), .B1(n12900), .Y(n8645)
         );
  NOR2X1 U7093 ( .A(n8648), .B(n8651), .Y(n8650) );
  INVX1 U7094 ( .A(n8652), .Y(n8651) );
  OAI21X1 U7095 ( .A0(n7857), .A1(n7607), .B0(n8653), .Y(n6863) );
  AOI22X1 U7096 ( .A0(n12902), .A1(n8654), .B0(n12901), .B1(n8655), .Y(n8653)
         );
  OAI21X1 U7097 ( .A0(n7857), .A1(n7634), .B0(n8656), .Y(n6862) );
  AOI22X1 U7098 ( .A0(n12903), .A1(n8654), .B0(n8655), .B1(n12902), .Y(n8656)
         );
  INVX1 U7099 ( .A(n8657), .Y(n6861) );
  AOI22X1 U7100 ( .A0(n8658), .A1(n7930), .B0(n12166), .B1(test_se), .Y(n8657)
         );
  MX2X1 U7101 ( .A(n8659), .B(n12489), .S0(n8660), .Y(n8658) );
  OAI21X1 U7102 ( .A0(n5899), .A1(n7857), .B0(n8661), .Y(n6860) );
  AOI22X1 U7103 ( .A0(n8662), .A1(n7930), .B0(n12771), .B1(n7909), .Y(n8661)
         );
  MX2X1 U7104 ( .A(n7258), .B(n12769), .S0(n12770), .Y(n8662) );
  OAI21X1 U7105 ( .A0(n5896), .A1(n7857), .B0(n8663), .Y(n6859) );
  AOI22X1 U7106 ( .A0(n7930), .A1(n8664), .B0(n12850), .B1(n7909), .Y(n8663)
         );
  OAI22X1 U7107 ( .A0(n12770), .A1(n7258), .B0(n8665), .B1(n7528), .Y(n8664)
         );
  AOI21X1 U7108 ( .A0(n8666), .A1(n8111), .B0(n12770), .Y(n8665) );
  NAND3X1 U7109 ( .A(n8659), .B(n7407), .C(n8667), .Y(n8666) );
  INVX1 U7110 ( .A(n8660), .Y(n8667) );
  NAND4X1 U7111 ( .A(n12931), .B(n12933), .C(g8719), .D(n7420), .Y(n8660) );
  NAND2X1 U7112 ( .A(n8668), .B(n8669), .Y(n8659) );
  NAND3X1 U7113 ( .A(n7244), .B(n7370), .C(n8670), .Y(n8669) );
  MX2X1 U7114 ( .A(n8671), .B(n8672), .S0(n7373), .Y(n8670) );
  AND2X1 U7115 ( .A(n7575), .B(n8673), .Y(n8672) );
  XOR2X1 U7116 ( .A(n12903), .B(n12902), .Y(n8673) );
  NOR2X1 U7117 ( .A(n12439), .B(n8674), .Y(n8671) );
  INVX1 U7118 ( .A(n8675), .Y(n8674) );
  XOR2X1 U7119 ( .A(n12415), .B(n12903), .Y(n8675) );
  OR2X1 U7120 ( .A(n8676), .B(n8677), .Y(n6858) );
  MX2X1 U7121 ( .A(test_se), .B(n8678), .S0(n7258), .Y(n8677) );
  NOR2X1 U7122 ( .A(n12769), .B(n7967), .Y(n8678) );
  AOI21X1 U7123 ( .A0(n7258), .A1(n7921), .B0(n7528), .Y(n8676) );
  NAND2X1 U7124 ( .A(n8679), .B(n8680), .Y(n6857) );
  MX2X1 U7125 ( .A(n12770), .B(n8681), .S0(n7847), .Y(n8680) );
  NAND2X1 U7126 ( .A(n8682), .B(n13035), .Y(n8681) );
  AOI22X1 U7127 ( .A0(n13034), .A1(n7908), .B0(n8683), .B1(n7930), .Y(n8679)
         );
  NOR2X1 U7128 ( .A(n13035), .B(n8682), .Y(n8683) );
  INVX1 U7129 ( .A(n8684), .Y(n8682) );
  NAND4X1 U7130 ( .A(n13045), .B(n13034), .C(n8476), .D(n7371), .Y(n8684) );
  NAND2X1 U7131 ( .A(n8685), .B(n8686), .Y(n6856) );
  AOI22X1 U7132 ( .A0(n8687), .A1(n13017), .B0(n8688), .B1(n8689), .Y(n8686)
         );
  NOR2X1 U7133 ( .A(n7494), .B(n8690), .Y(n8688) );
  AOI21X1 U7134 ( .A0(n8691), .A1(g7916), .B0(n7967), .Y(n8687) );
  AOI22X1 U7135 ( .A0(n13056), .A1(n7908), .B0(test_se), .B1(n7362), .Y(n8685)
         );
  INVX1 U7136 ( .A(n8692), .Y(n6855) );
  AOI22X1 U7137 ( .A0(n7930), .A1(n8693), .B0(n13017), .B1(test_se), .Y(n8692)
         );
  OAI21X1 U7138 ( .A0(n13071), .A1(n8694), .B0(n8695), .Y(n8693) );
  AOI22X1 U7139 ( .A0(n8696), .A1(n8697), .B0(n13068), .B1(n8698), .Y(n8695)
         );
  INVX1 U7140 ( .A(n8699), .Y(n8697) );
  AND2X1 U7141 ( .A(n8700), .B(n8701), .Y(n8696) );
  OAI21X1 U7142 ( .A0(n7857), .A1(n7609), .B0(n8702), .Y(n6854) );
  AOI22X1 U7143 ( .A0(n7930), .A1(n8703), .B0(n13061), .B1(n8704), .Y(n8702)
         );
  OAI21X1 U7144 ( .A0(test_se), .A1(n5888), .B0(n7919), .Y(n8704) );
  OAI21X1 U7145 ( .A0(n13061), .A1(n8705), .B0(g19334), .Y(n8703) );
  MX2X1 U7146 ( .A(n13042), .B(g13259), .S0(n7847), .Y(n6853) );
  OAI22X1 U7147 ( .A0(n7857), .A1(n7338), .B0(n8706), .B1(n7967), .Y(n6852) );
  AOI22X1 U7148 ( .A0(n8707), .A1(n8708), .B0(n12819), .B1(n8709), .Y(n8706)
         );
  NOR2X1 U7149 ( .A(n12818), .B(n12820), .Y(n8707) );
  MX2X1 U7150 ( .A(n12810), .B(n12799), .S0(n8710), .Y(n6851) );
  NAND2X1 U7151 ( .A(n8711), .B(n8712), .Y(n6850) );
  MX2X1 U7152 ( .A(n8713), .B(n8714), .S0(n7315), .Y(n8712) );
  NAND2X1 U7153 ( .A(n8715), .B(n7930), .Y(n8714) );
  AOI21X1 U7154 ( .A0(n8716), .A1(n8717), .B0(n7908), .Y(n8713) );
  NOR2X1 U7155 ( .A(n8718), .B(n8715), .Y(n8716) );
  NOR2X1 U7156 ( .A(n7515), .B(n8719), .Y(n8715) );
  AOI22X1 U7157 ( .A0(n12798), .A1(n8720), .B0(n12810), .B1(test_se), .Y(n8711) );
  OAI21X1 U7158 ( .A0(n8721), .A1(n7515), .B0(n8722), .Y(n6849) );
  AOI22X1 U7159 ( .A0(n8723), .A1(n8719), .B0(n8724), .B1(n7601), .Y(n8722) );
  OAI21X1 U7160 ( .A0(n8719), .A1(n7967), .B0(n8725), .Y(n8724) );
  INVX1 U7161 ( .A(n8720), .Y(n8725) );
  NOR2X1 U7162 ( .A(n8726), .B(n8727), .Y(n8723) );
  XOR2X1 U7163 ( .A(n12810), .B(n7515), .Y(n8726) );
  OAI21X1 U7164 ( .A0(n12797), .A1(n7930), .B0(n8728), .Y(n6848) );
  MX2X1 U7165 ( .A(n8729), .B(n8730), .S0(n7580), .Y(n8728) );
  NAND2X1 U7166 ( .A(n8731), .B(n8732), .Y(n8730) );
  MX2X1 U7167 ( .A(n12795), .B(n12796), .S0(n8710), .Y(n6847) );
  OAI21X1 U7168 ( .A0(n8710), .A1(n7240), .B0(n8733), .Y(n6846) );
  MX2X1 U7169 ( .A(n8734), .B(n8735), .S0(n12795), .Y(n8733) );
  AOI21X1 U7170 ( .A0(n8424), .A1(n12796), .B0(n8593), .Y(n8735) );
  NAND3X1 U7171 ( .A(n7930), .B(n7580), .C(n8424), .Y(n8734) );
  OAI21X1 U7172 ( .A0(n8710), .A1(n7307), .B0(n8736), .Y(n6845) );
  MX2X1 U7173 ( .A(n8737), .B(n7240), .S0(n7956), .Y(n8736) );
  NAND2X1 U7174 ( .A(n8424), .B(n7307), .Y(n8737) );
  INVX1 U7175 ( .A(n8738), .Y(n8710) );
  OAI22X1 U7176 ( .A0(n8729), .A1(n7651), .B0(n8739), .B1(n7307), .Y(n6844) );
  AOI21X1 U7177 ( .A0(n8731), .A1(n8740), .B0(n8593), .Y(n8739) );
  OAI21X1 U7178 ( .A0(n8729), .A1(n7215), .B0(n8741), .Y(n6843) );
  MX2X1 U7179 ( .A(n8742), .B(n8743), .S0(n7651), .Y(n8741) );
  NAND3X1 U7180 ( .A(n8732), .B(n7307), .C(n8731), .Y(n8743) );
  AOI21X1 U7181 ( .A0(n8744), .A1(n12794), .B0(n8593), .Y(n8742) );
  NOR2X1 U7182 ( .A(n8745), .B(n8746), .Y(n8744) );
  AOI21X1 U7183 ( .A0(n8746), .A1(n7930), .B0(n8720), .Y(n8729) );
  INVX1 U7184 ( .A(n8731), .Y(n8746) );
  OAI22X1 U7185 ( .A0(n7857), .A1(n7215), .B0(n8747), .B1(n7966), .Y(n6842) );
  AOI22X1 U7186 ( .A0(n8748), .A1(n8749), .B0(n12792), .B1(n8750), .Y(n8747)
         );
  NOR2X1 U7187 ( .A(n12791), .B(n12793), .Y(n8748) );
  MX2X1 U7188 ( .A(n12788), .B(n12776), .S0(n8751), .Y(n6841) );
  NAND2X1 U7189 ( .A(n8752), .B(n8753), .Y(n6840) );
  MX2X1 U7190 ( .A(n8754), .B(n8755), .S0(n7326), .Y(n8753) );
  NAND2X1 U7191 ( .A(n8756), .B(n7931), .Y(n8755) );
  AOI21X1 U7192 ( .A0(n8757), .A1(n8758), .B0(n7908), .Y(n8754) );
  NOR2X1 U7193 ( .A(test_se), .B(n8756), .Y(n8757) );
  NOR2X1 U7194 ( .A(n12775), .B(n8759), .Y(n8756) );
  AOI22X1 U7195 ( .A0(n8760), .A1(n7432), .B0(n12788), .B1(test_se), .Y(n8752)
         );
  OAI21X1 U7196 ( .A0(n12775), .A1(n8721), .B0(n8761), .Y(n6839) );
  AOI22X1 U7197 ( .A0(n8762), .A1(n8763), .B0(n12774), .B1(n8764), .Y(n8761)
         );
  OAI21X1 U7198 ( .A0(n8759), .A1(n7966), .B0(n8765), .Y(n8764) );
  XOR2X1 U7199 ( .A(n12788), .B(n7432), .Y(n8763) );
  AND2X1 U7200 ( .A(n8766), .B(n8759), .Y(n8762) );
  OAI21X1 U7201 ( .A0(n7856), .A1(n7784), .B0(n8767), .Y(n6838) );
  AOI21X1 U7202 ( .A0(n7908), .A1(g20652), .B0(n8768), .Y(n8767) );
  AOI21X1 U7203 ( .A0(n8769), .A1(n7741), .B0(n7966), .Y(n8768) );
  OAI21X1 U7204 ( .A0(n7856), .A1(n7785), .B0(n8770), .Y(n6837) );
  AOI22X1 U7205 ( .A0(n7931), .A1(n8771), .B0(n12681), .B1(n7908), .Y(n8770)
         );
  NAND4X1 U7206 ( .A(n8772), .B(n8773), .C(n7744), .D(n7318), .Y(n8771) );
  AOI21X1 U7207 ( .A0(test_se), .A1(n7786), .B0(n8774), .Y(n6836) );
  OAI21X1 U7208 ( .A0(n12671), .A1(n7921), .B0(n8775), .Y(n8774) );
  NAND3X1 U7209 ( .A(n7931), .B(n7742), .C(n8776), .Y(n8775) );
  OAI21X1 U7210 ( .A0(n7856), .A1(n7742), .B0(n8777), .Y(n6835) );
  AOI22X1 U7211 ( .A0(n7931), .A1(n8778), .B0(n12659), .B1(n7908), .Y(n8777)
         );
  NAND3X1 U7212 ( .A(n7343), .B(n7670), .C(n8779), .Y(n8778) );
  OAI21X1 U7213 ( .A0(n7856), .A1(n7670), .B0(n8780), .Y(n6834) );
  AOI22X1 U7214 ( .A0(n12657), .A1(n7908), .B0(n12658), .B1(n7931), .Y(n8780)
         );
  MX2X1 U7215 ( .A(n12656), .B(n12658), .S0(n7956), .Y(n6833) );
  OAI21X1 U7216 ( .A0(n7856), .A1(n7706), .B0(n8781), .Y(n6832) );
  AOI22X1 U7217 ( .A0(n7931), .A1(n8782), .B0(n12660), .B1(n7908), .Y(n8781)
         );
  NAND3X1 U7218 ( .A(n8783), .B(n7671), .C(n8784), .Y(n8782) );
  OAI21X1 U7219 ( .A0(n7856), .A1(n7671), .B0(n8785), .Y(n6831) );
  AOI22X1 U7220 ( .A0(n12656), .A1(n7908), .B0(n12654), .B1(n7931), .Y(n8785)
         );
  OR2X1 U7221 ( .A(n8786), .B(n7931), .Y(n6830) );
  MX2X1 U7222 ( .A(n12654), .B(n12655), .S0(n7847), .Y(n8786) );
  OAI21X1 U7223 ( .A0(n7856), .A1(n7834), .B0(n8787), .Y(n6829) );
  AOI22X1 U7224 ( .A0(n12654), .A1(n7908), .B0(n12651), .B1(n7931), .Y(n8787)
         );
  OAI21X1 U7225 ( .A0(n7856), .A1(n7707), .B0(n8788), .Y(n6828) );
  AOI22X1 U7226 ( .A0(n7931), .A1(n8789), .B0(n7908), .B1(n12652), .Y(n8788)
         );
  NAND3X1 U7227 ( .A(n7231), .B(n7672), .C(n7339), .Y(n8789) );
  OAI21X1 U7228 ( .A0(n7856), .A1(n7672), .B0(n8790), .Y(n6827) );
  MX2X1 U7229 ( .A(n8791), .B(n8792), .S0(n7539), .Y(n8790) );
  OR2X1 U7230 ( .A(n7966), .B(n5856), .Y(n8792) );
  AOI21X1 U7231 ( .A0(n5856), .A1(n7856), .B0(n7907), .Y(n8791) );
  OAI21X1 U7232 ( .A0(n12663), .A1(n7856), .B0(n8793), .Y(n6826) );
  AOI22X1 U7233 ( .A0(n12651), .A1(n7907), .B0(n12646), .B1(n7931), .Y(n8793)
         );
  OAI21X1 U7234 ( .A0(n7855), .A1(n7708), .B0(n8794), .Y(n6825) );
  AOI22X1 U7235 ( .A0(n7931), .A1(n8795), .B0(n12647), .B1(n7907), .Y(n8794)
         );
  OR2X1 U7236 ( .A(n8796), .B(n8797), .Y(n8795) );
  NAND3X1 U7237 ( .A(n8798), .B(n8776), .C(n12663), .Y(n8797) );
  INVX1 U7238 ( .A(n8799), .Y(n8776) );
  NAND4X1 U7239 ( .A(n8800), .B(n8801), .C(n8802), .D(n8803), .Y(n8799) );
  NAND4X1 U7240 ( .A(n8772), .B(n8769), .C(n8280), .D(n7673), .Y(n8796) );
  NOR2X1 U7241 ( .A(n8804), .B(n8805), .Y(n8280) );
  NOR2X1 U7242 ( .A(n8806), .B(n8807), .Y(n8769) );
  OAI21X1 U7243 ( .A0(n7855), .A1(n7673), .B0(n8808), .Y(n6824) );
  AOI22X1 U7244 ( .A0(n12646), .A1(n7907), .B0(n12644), .B1(n7931), .Y(n8808)
         );
  OR2X1 U7245 ( .A(n8809), .B(n7931), .Y(n6823) );
  MX2X1 U7246 ( .A(n12644), .B(n12645), .S0(n7848), .Y(n8809) );
  OAI21X1 U7247 ( .A0(n7856), .A1(n7787), .B0(n8810), .Y(n6822) );
  AOI22X1 U7248 ( .A0(n12644), .A1(n7907), .B0(n12659), .B1(n7931), .Y(n8810)
         );
  OAI21X1 U7249 ( .A0(n7855), .A1(n7709), .B0(n8811), .Y(n6821) );
  AOI22X1 U7250 ( .A0(n7931), .A1(n8812), .B0(n12643), .B1(n7907), .Y(n8811)
         );
  NAND3X1 U7251 ( .A(n13017), .B(n7674), .C(n12965), .Y(n8812) );
  OAI21X1 U7252 ( .A0(n7855), .A1(n7674), .B0(n8813), .Y(n6820) );
  AOI21X1 U7253 ( .A0(n12662), .A1(n7907), .B0(n8814), .Y(n8813) );
  AOI21X1 U7254 ( .A0(n7352), .A1(n7835), .B0(n7966), .Y(n8814) );
  OAI21X1 U7255 ( .A0(n7855), .A1(n7743), .B0(n8815), .Y(n6819) );
  AOI21X1 U7256 ( .A0(n12640), .A1(n7907), .B0(n8163), .Y(n8815) );
  OAI21X1 U7257 ( .A0(n7855), .A1(n7744), .B0(n8816), .Y(n6818) );
  AOI22X1 U7258 ( .A0(n12668), .A1(n7907), .B0(n12669), .B1(n7931), .Y(n8816)
         );
  INVX1 U7259 ( .A(n8817), .Y(n6817) );
  AOI22X1 U7260 ( .A0(n12669), .A1(n8593), .B0(n12667), .B1(n7931), .Y(n8817)
         );
  INVX1 U7261 ( .A(n8818), .Y(n6816) );
  AOI22X1 U7262 ( .A0(n12642), .A1(n7907), .B0(n12639), .B1(test_se), .Y(n8818) );
  OAI21X1 U7263 ( .A0(n489), .A1(n7855), .B0(n8819), .Y(n6815) );
  AOI21X1 U7264 ( .A0(n12638), .A1(n7907), .B0(n8820), .Y(n8819) );
  NAND2X1 U7265 ( .A(n8821), .B(n8822), .Y(n6814) );
  MX2X1 U7266 ( .A(n8823), .B(n8824), .S0(n12602), .Y(n8822) );
  INVX1 U7267 ( .A(n8825), .Y(n8824) );
  OAI21X1 U7268 ( .A0(n8826), .A1(n8827), .B0(n7923), .Y(n8823) );
  XOR2X1 U7269 ( .A(n8828), .B(n8829), .Y(n8827) );
  AOI22X1 U7270 ( .A0(n12634), .A1(n7907), .B0(n12637), .B1(test_se), .Y(n8821) );
  OAI21X1 U7271 ( .A0(n8830), .A1(n7229), .B0(n8831), .Y(n6813) );
  NOR2X1 U7272 ( .A(n8832), .B(n8833), .Y(n8831) );
  AOI21X1 U7273 ( .A0(n7921), .A1(n8834), .B0(n12602), .Y(n8833) );
  NAND3X1 U7274 ( .A(n7675), .B(n7855), .C(n8835), .Y(n8834) );
  AOI21X1 U7275 ( .A0(n7855), .A1(n8836), .B0(n7675), .Y(n8832) );
  NAND3X1 U7276 ( .A(n12602), .B(g35), .C(n8835), .Y(n8836) );
  OAI21X1 U7277 ( .A0(n8837), .A1(n7558), .B0(n8838), .Y(n6812) );
  MX2X1 U7278 ( .A(n8839), .B(n7229), .S0(n7956), .Y(n8838) );
  NAND2X1 U7279 ( .A(n8510), .B(n7558), .Y(n8839) );
  OAI21X1 U7280 ( .A0(n12597), .A1(n8830), .B0(n8840), .Y(n6811) );
  OAI21X1 U7281 ( .A0(n8835), .A1(n8593), .B0(n12598), .Y(n8840) );
  OAI21X1 U7282 ( .A0(n12689), .A1(n8830), .B0(n8841), .Y(n6810) );
  MX2X1 U7283 ( .A(n8842), .B(n8843), .S0(n12597), .Y(n8841) );
  NAND3X1 U7284 ( .A(n7931), .B(n7558), .C(n8835), .Y(n8843) );
  AOI21X1 U7285 ( .A0(n12598), .A1(n8835), .B0(n8593), .Y(n8842) );
  OAI21X1 U7286 ( .A0(n8830), .A1(n7559), .B0(n8844), .Y(n6809) );
  MX2X1 U7287 ( .A(n8845), .B(n12689), .S0(n7955), .Y(n8844) );
  NAND2X1 U7288 ( .A(n8835), .B(n7559), .Y(n8845) );
  OR2X1 U7289 ( .A(n7966), .B(n8835), .Y(n8830) );
  NOR2X1 U7290 ( .A(n8846), .B(n8826), .Y(n8835) );
  MX2X1 U7291 ( .A(n12595), .B(n12596), .S0(n8837), .Y(n6808) );
  OAI21X1 U7292 ( .A0(n8837), .A1(n7644), .B0(n8847), .Y(n6807) );
  MX2X1 U7293 ( .A(n8848), .B(n8849), .S0(n12595), .Y(n8847) );
  AOI21X1 U7294 ( .A0(n12596), .A1(n8510), .B0(n8593), .Y(n8849) );
  NAND3X1 U7295 ( .A(n7931), .B(n7559), .C(n8510), .Y(n8848) );
  INVX1 U7296 ( .A(n8508), .Y(n8837) );
  OAI21X1 U7297 ( .A0(n7855), .A1(n7745), .B0(n8850), .Y(n6806) );
  NAND3X1 U7298 ( .A(n7217), .B(n7301), .C(n7931), .Y(n8850) );
  NAND2X1 U7299 ( .A(n8851), .B(n8852), .Y(n6805) );
  MX2X1 U7300 ( .A(n8853), .B(n7301), .S0(n7955), .Y(n8851) );
  OAI22X1 U7301 ( .A0(n8854), .A1(n12600), .B0(n7564), .B1(n7931), .Y(n6804)
         );
  XOR2X1 U7302 ( .A(n7217), .B(n8855), .Y(n6803) );
  NAND2X1 U7303 ( .A(n12601), .B(n7931), .Y(n8855) );
  MX2X1 U7304 ( .A(n8856), .B(n12601), .S0(n7955), .Y(n6802) );
  NAND3X1 U7305 ( .A(n8857), .B(n8858), .C(n8859), .Y(n8856) );
  NAND2X1 U7306 ( .A(n12636), .B(n7217), .Y(n8859) );
  INVX1 U7307 ( .A(n8860), .Y(n6801) );
  AOI22X1 U7308 ( .A0(n12636), .A1(n7932), .B0(n12638), .B1(test_se), .Y(n8860) );
  OAI21X1 U7309 ( .A0(n8534), .A1(n8861), .B0(n8862), .Y(n6800) );
  MX2X1 U7310 ( .A(n8863), .B(n7480), .S0(n7955), .Y(n8862) );
  NAND2X1 U7311 ( .A(n12616), .B(n8861), .Y(n8863) );
  OR2X1 U7312 ( .A(n8864), .B(n8865), .Y(n8861) );
  NAND2X1 U7313 ( .A(n8866), .B(n8867), .Y(n6799) );
  MX2X1 U7314 ( .A(n8868), .B(n8534), .S0(n8869), .Y(n8867) );
  NOR2X1 U7315 ( .A(n8864), .B(n8852), .Y(n8869) );
  NAND2X1 U7316 ( .A(n12615), .B(n7932), .Y(n8868) );
  AOI22X1 U7317 ( .A0(n12616), .A1(n7906), .B0(n12631), .B1(test_se), .Y(n8866) );
  NAND2X1 U7318 ( .A(n8870), .B(n8871), .Y(n6798) );
  MX2X1 U7319 ( .A(n8872), .B(n8534), .S0(n8873), .Y(n8871) );
  NOR2X1 U7320 ( .A(n8853), .B(n8864), .Y(n8873) );
  NAND2X1 U7321 ( .A(n12613), .B(n7932), .Y(n8872) );
  AOI22X1 U7322 ( .A0(n12615), .A1(n7906), .B0(n12623), .B1(test_se), .Y(n8870) );
  NAND2X1 U7323 ( .A(n8874), .B(n8875), .Y(n6797) );
  MX2X1 U7324 ( .A(n8876), .B(n8534), .S0(n8877), .Y(n8875) );
  NOR2X1 U7325 ( .A(n8854), .B(n8864), .Y(n8877) );
  NAND2X1 U7326 ( .A(n7932), .B(n7225), .Y(n8876) );
  AOI22X1 U7327 ( .A0(n12613), .A1(n7906), .B0(n12622), .B1(test_se), .Y(n8874) );
  NAND2X1 U7328 ( .A(n8878), .B(n8879), .Y(n6796) );
  MX2X1 U7329 ( .A(n8880), .B(n8534), .S0(n8881), .Y(n8879) );
  NOR2X1 U7330 ( .A(n8854), .B(n8882), .Y(n8881) );
  NAND2X1 U7331 ( .A(n12626), .B(n7932), .Y(n8880) );
  AOI22X1 U7332 ( .A0(n12625), .A1(n7906), .B0(test_se), .B1(n7225), .Y(n8878)
         );
  NAND2X1 U7333 ( .A(n8883), .B(n8884), .Y(n6795) );
  MX2X1 U7334 ( .A(n8885), .B(n8534), .S0(n8886), .Y(n8884) );
  NOR2X1 U7335 ( .A(n8854), .B(n8858), .Y(n8886) );
  NAND2X1 U7336 ( .A(n12620), .B(n7932), .Y(n8885) );
  AOI22X1 U7337 ( .A0(n12628), .A1(n7906), .B0(n12626), .B1(test_se), .Y(n8883) );
  NAND2X1 U7338 ( .A(n8887), .B(n8888), .Y(n6794) );
  MX2X1 U7339 ( .A(n8889), .B(n8534), .S0(n8890), .Y(n8888) );
  NOR2X1 U7340 ( .A(n8891), .B(n8854), .Y(n8890) );
  NAND2X1 U7341 ( .A(n12591), .B(n12592), .Y(n8854) );
  NAND2X1 U7342 ( .A(n12621), .B(n7932), .Y(n8889) );
  AOI22X1 U7343 ( .A0(n12622), .A1(n7906), .B0(n12620), .B1(test_se), .Y(n8887) );
  OAI21X1 U7344 ( .A0(n7932), .A1(n7788), .B0(n8892), .Y(n6793) );
  AOI22X1 U7345 ( .A0(n12614), .A1(n8508), .B0(n8893), .B1(n8510), .Y(n8892)
         );
  NOR2X1 U7346 ( .A(n7966), .B(n8510), .Y(n8508) );
  NOR2X1 U7347 ( .A(n7217), .B(n8891), .Y(n8510) );
  NAND2X1 U7348 ( .A(n8894), .B(n8895), .Y(n6792) );
  AOI21X1 U7349 ( .A0(n12587), .A1(n8896), .B0(n8825), .Y(n8895) );
  NOR2X1 U7350 ( .A(n8897), .B(n8829), .Y(n8825) );
  AOI21X1 U7351 ( .A0(n12614), .A1(n8828), .B0(n8898), .Y(n8829) );
  MX2X1 U7352 ( .A(n8899), .B(n8900), .S0(n7422), .Y(n8898) );
  NAND4X1 U7353 ( .A(n8901), .B(n8902), .C(n8903), .D(n8904), .Y(n8900) );
  NAND3X1 U7354 ( .A(n8905), .B(g16874), .C(n12618), .Y(n8904) );
  NAND2X1 U7355 ( .A(n8906), .B(n8907), .Y(n8903) );
  INVX1 U7356 ( .A(n8908), .Y(n8906) );
  AOI22X1 U7357 ( .A0(n12620), .A1(g16686), .B0(n12619), .B1(g16624), .Y(n8908) );
  OR2X1 U7358 ( .A(n12632), .B(n8909), .Y(n8902) );
  MX2X1 U7359 ( .A(n8910), .B(n8911), .S0(n7361), .Y(n8909) );
  NAND2X1 U7360 ( .A(n12628), .B(g13865), .Y(n8911) );
  AOI22X1 U7361 ( .A0(n12629), .A1(g14421), .B0(n12631), .B1(n12630), .Y(n8910) );
  MX2X1 U7362 ( .A(n8912), .B(n8913), .S0(g11349), .Y(n8901) );
  AOI21X1 U7363 ( .A0(n12624), .A1(n8905), .B0(n8914), .Y(n8913) );
  INVX1 U7364 ( .A(n8915), .Y(n8912) );
  NAND4X1 U7365 ( .A(n8916), .B(n8917), .C(n8918), .D(n8919), .Y(n8899) );
  NAND3X1 U7366 ( .A(n8920), .B(g13865), .C(n12613), .Y(n8919) );
  NAND3X1 U7367 ( .A(g16686), .B(n7225), .C(n8905), .Y(n8918) );
  OR2X1 U7368 ( .A(n12633), .B(n8921), .Y(n8917) );
  MX2X1 U7369 ( .A(n8922), .B(n8923), .S0(n7242), .Y(n8921) );
  AOI22X1 U7370 ( .A0(n12616), .A1(g14421), .B0(n12617), .B1(n12630), .Y(n8923) );
  AOI22X1 U7371 ( .A0(n12615), .A1(g16874), .B0(g11349), .B1(n7278), .Y(n8922)
         );
  INVX1 U7372 ( .A(n8924), .Y(n8916) );
  MX2X1 U7373 ( .A(n8914), .B(n8915), .S0(g11349), .Y(n8924) );
  NAND3X1 U7374 ( .A(n8925), .B(n8926), .C(n8927), .Y(n8915) );
  NAND3X1 U7375 ( .A(n8905), .B(g16718), .C(n12625), .Y(n8927) );
  NAND3X1 U7376 ( .A(n8928), .B(g16603), .C(n12626), .Y(n8926) );
  NAND3X1 U7377 ( .A(n8920), .B(g13895), .C(n12627), .Y(n8925) );
  NAND3X1 U7378 ( .A(n8929), .B(n8930), .C(n8931), .Y(n8914) );
  NAND3X1 U7379 ( .A(n8920), .B(g16603), .C(n12621), .Y(n8931) );
  NAND3X1 U7380 ( .A(n8928), .B(g13895), .C(n12623), .Y(n8930) );
  NAND3X1 U7381 ( .A(n8907), .B(g16718), .C(n12622), .Y(n8929) );
  INVX1 U7382 ( .A(n8846), .Y(n8828) );
  NAND3X1 U7383 ( .A(n12635), .B(g16624), .C(n8905), .Y(n8846) );
  AOI22X1 U7384 ( .A0(n12614), .A1(n7906), .B0(n12630), .B1(test_se), .Y(n8894) );
  NAND2X1 U7385 ( .A(n8932), .B(n8933), .Y(n6791) );
  MX2X1 U7386 ( .A(n8934), .B(n8935), .S0(n8936), .Y(n8933) );
  NAND2X1 U7387 ( .A(n7932), .B(n7422), .Y(n8934) );
  AOI22X1 U7388 ( .A0(n12630), .A1(n7906), .B0(n12587), .B1(test_se), .Y(n8932) );
  NOR2X1 U7389 ( .A(n8937), .B(n8938), .Y(n6790) );
  MX2X1 U7390 ( .A(n12586), .B(n7422), .S0(n7948), .Y(n8938) );
  NOR2X1 U7391 ( .A(n8937), .B(n7652), .Y(n6789) );
  NOR2X1 U7392 ( .A(n8935), .B(n8936), .Y(n8937) );
  NAND4X1 U7393 ( .A(g16718), .B(g16603), .C(g13895), .D(g11349), .Y(n8936) );
  INVX1 U7394 ( .A(n8820), .Y(n8935) );
  NOR2X1 U7395 ( .A(n7422), .B(n7966), .Y(n8820) );
  OAI21X1 U7396 ( .A0(n12604), .A1(n7855), .B0(n8939), .Y(n6788) );
  AOI22X1 U7397 ( .A0(n8940), .A1(n8941), .B0(n12302), .B1(n8942), .Y(n8939)
         );
  OAI21X1 U7398 ( .A0(n7966), .A1(n8943), .B0(n8944), .Y(n8942) );
  AOI21X1 U7399 ( .A0(n8945), .A1(n8946), .B0(n8897), .Y(n8940) );
  INVX1 U7400 ( .A(n8947), .Y(n8946) );
  MX2X1 U7401 ( .A(n8920), .B(n8928), .S0(n7652), .Y(n8947) );
  NOR2X1 U7402 ( .A(n12633), .B(n12632), .Y(n8928) );
  NOR2X1 U7403 ( .A(n7361), .B(n12632), .Y(n8920) );
  INVX1 U7404 ( .A(n8948), .Y(n8945) );
  MX2X1 U7405 ( .A(n8905), .B(n8907), .S0(n7624), .Y(n8948) );
  NOR2X1 U7406 ( .A(n7242), .B(n12633), .Y(n8907) );
  NOR2X1 U7407 ( .A(n7361), .B(n7242), .Y(n8905) );
  OAI21X1 U7408 ( .A0(n7855), .A1(n7789), .B0(n8949), .Y(n6787) );
  AOI21X1 U7409 ( .A0(n8950), .A1(n7363), .B0(n8951), .Y(n8949) );
  AOI21X1 U7410 ( .A0(n7921), .A1(n8952), .B0(n12608), .Y(n8951) );
  NAND3X1 U7411 ( .A(n8953), .B(n7855), .C(n8954), .Y(n8952) );
  OAI21X1 U7412 ( .A0(n12610), .A1(n7932), .B0(n8955), .Y(n6786) );
  MX2X1 U7413 ( .A(n8953), .B(n8956), .S0(n7247), .Y(n8955) );
  NAND2X1 U7414 ( .A(n8957), .B(n8958), .Y(n6785) );
  AOI22X1 U7415 ( .A0(n8950), .A1(n7379), .B0(n8523), .B1(n7932), .Y(n8958) );
  AOI21X1 U7416 ( .A0(n7906), .A1(n7247), .B0(n8959), .Y(n8957) );
  MX2X1 U7417 ( .A(n12306), .B(n8960), .S0(n7849), .Y(n8959) );
  NOR2X1 U7418 ( .A(n8616), .B(n8953), .Y(n8960) );
  INVX1 U7419 ( .A(n8579), .Y(n8616) );
  INVX1 U7420 ( .A(n8961), .Y(n6784) );
  AOI22X1 U7421 ( .A0(n12390), .A1(n7932), .B0(test_se), .B1(n7379), .Y(n8961)
         );
  INVX1 U7422 ( .A(n8962), .Y(n6783) );
  AOI22X1 U7423 ( .A0(n12390), .A1(n8593), .B0(n12389), .B1(n7932), .Y(n8962)
         );
  INVX1 U7424 ( .A(n8963), .Y(n6782) );
  AOI22X1 U7425 ( .A0(n12389), .A1(n8593), .B0(n12388), .B1(n7932), .Y(n8963)
         );
  OAI21X1 U7426 ( .A0(n7855), .A1(n7746), .B0(n8964), .Y(n6781) );
  AOI22X1 U7427 ( .A0(n8965), .A1(n7932), .B0(n12302), .B1(n8966), .Y(n8964)
         );
  OAI21X1 U7428 ( .A0(test_se), .A1(n8943), .B0(n7919), .Y(n8966) );
  NOR2X1 U7429 ( .A(n12604), .B(n8941), .Y(n8965) );
  INVX1 U7430 ( .A(n8943), .Y(n8941) );
  NAND2X1 U7431 ( .A(n8339), .B(n8615), .Y(n8943) );
  INVX1 U7432 ( .A(n8603), .Y(n8339) );
  NAND3X1 U7433 ( .A(n7363), .B(n7250), .C(n12608), .Y(n8603) );
  OAI21X1 U7434 ( .A0(n7855), .A1(n7836), .B0(n8967), .Y(n6780) );
  AOI22X1 U7435 ( .A0(n8968), .A1(n7932), .B0(n7906), .B1(n7228), .Y(n8967) );
  NOR2X1 U7436 ( .A(n12427), .B(n12449), .Y(n8968) );
  OAI21X1 U7437 ( .A0(n7854), .A1(n7685), .B0(n8969), .Y(n6779) );
  AOI22X1 U7438 ( .A0(n8970), .A1(n8971), .B0(n7906), .B1(n7364), .Y(n8969) );
  XOR2X1 U7439 ( .A(n8972), .B(n7359), .Y(n8970) );
  OAI21X1 U7440 ( .A0(n12446), .A1(n7932), .B0(n8973), .Y(n6778) );
  MX2X1 U7441 ( .A(n8974), .B(n8975), .S0(n7355), .Y(n8973) );
  NAND2X1 U7442 ( .A(n8971), .B(n8976), .Y(n8975) );
  NAND2X1 U7443 ( .A(n8977), .B(n12444), .Y(n8974) );
  INVX1 U7444 ( .A(n8978), .Y(n6777) );
  AOI22X1 U7445 ( .A0(n8979), .A1(n8971), .B0(n7966), .B1(n7355), .Y(n8978) );
  XOR2X1 U7446 ( .A(n8980), .B(n7410), .Y(n8979) );
  OAI21X1 U7447 ( .A0(n12443), .A1(n8721), .B0(n8981), .Y(n6776) );
  MX2X1 U7448 ( .A(n8982), .B(n8983), .S0(n12445), .Y(n8981) );
  NAND2X1 U7449 ( .A(n8984), .B(n12444), .Y(n8983) );
  NAND2X1 U7450 ( .A(n8971), .B(n8985), .Y(n8982) );
  INVX1 U7451 ( .A(n8986), .Y(n8971) );
  OAI22X1 U7452 ( .A0(n12444), .A1(n8986), .B0(n12445), .B1(n8987), .Y(n6775)
         );
  AOI21X1 U7453 ( .A0(n8984), .A1(n12444), .B0(n7966), .Y(n8987) );
  INVX1 U7454 ( .A(n8985), .Y(n8984) );
  NAND2X1 U7455 ( .A(n8980), .B(n7410), .Y(n8985) );
  NOR2X1 U7456 ( .A(n8976), .B(n12442), .Y(n8980) );
  OAI21X1 U7457 ( .A0(n12444), .A1(n8976), .B0(n7923), .Y(n8986) );
  INVX1 U7458 ( .A(n8977), .Y(n8976) );
  NOR2X1 U7459 ( .A(n8988), .B(n12446), .Y(n8977) );
  OAI21X1 U7460 ( .A0(n12444), .A1(n7854), .B0(n8989), .Y(n6774) );
  MX2X1 U7461 ( .A(n8990), .B(n8991), .S0(n12456), .Y(n8989) );
  NAND2X1 U7462 ( .A(n8992), .B(n7413), .Y(n8991) );
  AOI21X1 U7463 ( .A0(n8993), .A1(n12455), .B0(n7906), .Y(n8990) );
  NOR2X1 U7464 ( .A(test_se), .B(n7245), .Y(n8993) );
  OAI21X1 U7465 ( .A0(n12455), .A1(n7932), .B0(n8994), .Y(n6773) );
  MX2X1 U7466 ( .A(n8995), .B(n8996), .S0(n7277), .Y(n8994) );
  NAND2X1 U7467 ( .A(n8992), .B(n8997), .Y(n8996) );
  INVX1 U7468 ( .A(n8998), .Y(n8997) );
  NAND2X1 U7469 ( .A(n8998), .B(n12450), .Y(n8995) );
  OAI21X1 U7470 ( .A0(n12454), .A1(n8721), .B0(n8999), .Y(n6772) );
  MX2X1 U7471 ( .A(n9000), .B(n9001), .S0(n7276), .Y(n8999) );
  NAND2X1 U7472 ( .A(n8992), .B(n9002), .Y(n9001) );
  OR2X1 U7473 ( .A(n9002), .B(n7245), .Y(n9000) );
  NAND2X1 U7474 ( .A(n8998), .B(n7277), .Y(n9002) );
  NOR2X1 U7475 ( .A(n12456), .B(n12455), .Y(n8998) );
  OAI21X1 U7476 ( .A0(n12385), .A1(n7921), .B0(n9003), .Y(n6771) );
  MX2X1 U7477 ( .A(n12456), .B(n9004), .S0(n7850), .Y(n9003) );
  NAND2X1 U7478 ( .A(n12450), .B(n8139), .Y(n9004) );
  INVX1 U7479 ( .A(n9005), .Y(n8139) );
  NAND3X1 U7480 ( .A(n7413), .B(n7276), .C(n12456), .Y(n9005) );
  INVX1 U7481 ( .A(n9006), .Y(n6770) );
  AOI22X1 U7482 ( .A0(n8992), .A1(n12456), .B0(test_se), .B1(n7276), .Y(n9006)
         );
  NOR2X1 U7483 ( .A(n7245), .B(n7966), .Y(n8992) );
  INVX1 U7484 ( .A(n9007), .Y(n6769) );
  AOI22X1 U7485 ( .A0(n9008), .A1(n9009), .B0(test_se), .B1(n7245), .Y(n9007)
         );
  INVX1 U7486 ( .A(n8625), .Y(n9009) );
  NAND3X1 U7487 ( .A(n12404), .B(n7608), .C(n12403), .Y(n8625) );
  OAI21X1 U7488 ( .A0(n7854), .A1(n7608), .B0(n9010), .Y(n6768) );
  MX2X1 U7489 ( .A(n9011), .B(n9012), .S0(n7360), .Y(n9010) );
  AOI21X1 U7490 ( .A0(n7577), .A1(n7855), .B0(n7905), .Y(n9012) );
  NAND2X1 U7491 ( .A(n9008), .B(n12999), .Y(n9011) );
  OAI21X1 U7492 ( .A0(n7932), .A1(n7577), .B0(n9013), .Y(n6767) );
  MX2X1 U7493 ( .A(n9014), .B(n9015), .S0(n7433), .Y(n9013) );
  NAND2X1 U7494 ( .A(n9008), .B(n9014), .Y(n9015) );
  NOR2X1 U7495 ( .A(n7966), .B(n9016), .Y(n9008) );
  MX2X1 U7496 ( .A(n9017), .B(n7433), .S0(n7954), .Y(n6766) );
  MX2X1 U7497 ( .A(n9018), .B(n9019), .S0(n7653), .Y(n9017) );
  NOR2X1 U7498 ( .A(n12998), .B(n9018), .Y(n9019) );
  OAI21X1 U7499 ( .A0(n9020), .A1(n7653), .B0(n9021), .Y(n6765) );
  NAND3X1 U7500 ( .A(n7932), .B(n9018), .C(n12998), .Y(n9021) );
  AOI21X1 U7501 ( .A0(n9022), .A1(n7546), .B0(n8593), .Y(n9020) );
  MX2X1 U7502 ( .A(n12998), .B(n12995), .S0(n7850), .Y(n6764) );
  OAI21X1 U7503 ( .A0(n7854), .A1(n7747), .B0(n9023), .Y(n6762) );
  AOI22X1 U7504 ( .A0(n7932), .A1(n9024), .B0(n12238), .B1(n7905), .Y(n9023)
         );
  OAI21X1 U7505 ( .A0(n8359), .A1(n9025), .B0(n9026), .Y(n9024) );
  MX2X1 U7506 ( .A(n9027), .B(n12239), .S0(n9028), .Y(n9026) );
  NAND2X1 U7507 ( .A(n8359), .B(n9025), .Y(n9027) );
  NAND2X1 U7508 ( .A(n9029), .B(n7578), .Y(n9025) );
  MX2X1 U7509 ( .A(n9030), .B(n9031), .S0(n7415), .Y(n8359) );
  NAND4X1 U7510 ( .A(n9032), .B(n9033), .C(n9034), .D(n9035), .Y(n9031) );
  OR2X1 U7511 ( .A(n9036), .B(n9037), .Y(n9035) );
  AOI22X1 U7512 ( .A0(n12352), .A1(g13049), .B0(n12353), .B1(n12367), .Y(n9036) );
  AOI22X1 U7513 ( .A0(n9038), .A1(n12355), .B0(n9039), .B1(n12354), .Y(n9034)
         );
  NOR2X1 U7514 ( .A(n5258), .B(n9040), .Y(n9039) );
  NOR2X1 U7515 ( .A(n5259), .B(n9041), .Y(n9038) );
  OR2X1 U7516 ( .A(n9042), .B(n9043), .Y(n9033) );
  AOI22X1 U7517 ( .A0(g17678), .A1(n7226), .B0(n12371), .B1(g17604), .Y(n9042)
         );
  MX2X1 U7518 ( .A(n9044), .B(n9045), .S0(g12300), .Y(n9032) );
  AOI21X1 U7519 ( .A0(n9046), .A1(n7440), .B0(n9047), .Y(n9045) );
  INVX1 U7520 ( .A(n9048), .Y(n9044) );
  NAND4X1 U7521 ( .A(n9049), .B(n9050), .C(n9051), .D(n9052), .Y(n9030) );
  OR2X1 U7522 ( .A(n9053), .B(n9041), .Y(n9052) );
  AOI22X1 U7523 ( .A0(n12358), .A1(g17678), .B0(n12357), .B1(g17604), .Y(n9053) );
  AOI22X1 U7524 ( .A0(n9054), .A1(n12369), .B0(n9055), .B1(n12370), .Y(n9051)
         );
  NOR2X1 U7525 ( .A(n5259), .B(n9043), .Y(n9055) );
  INVX1 U7526 ( .A(n9056), .Y(n9043) );
  NOR2X1 U7527 ( .A(n5258), .B(n9037), .Y(n9054) );
  INVX1 U7528 ( .A(n9057), .Y(n9037) );
  OR2X1 U7529 ( .A(n9058), .B(n9040), .Y(n9050) );
  INVX1 U7530 ( .A(n9059), .Y(n9040) );
  AOI22X1 U7531 ( .A0(n12366), .A1(g13049), .B0(n12367), .B1(n12368), .Y(n9058) );
  MX2X1 U7532 ( .A(n9060), .B(n9061), .S0(g12300), .Y(n9049) );
  AOI21X1 U7533 ( .A0(n12362), .A1(n9056), .B0(n9048), .Y(n9061) );
  NAND3X1 U7534 ( .A(n9062), .B(n9063), .C(n9064), .Y(n9048) );
  NAND3X1 U7535 ( .A(n9059), .B(g17580), .C(n12360), .Y(n9064) );
  NAND3X1 U7536 ( .A(n9046), .B(g17711), .C(n12361), .Y(n9063) );
  NAND3X1 U7537 ( .A(n9057), .B(g14694), .C(n12359), .Y(n9062) );
  INVX1 U7538 ( .A(n9047), .Y(n9060) );
  NAND3X1 U7539 ( .A(n9065), .B(n9066), .C(n9067), .Y(n9047) );
  NAND3X1 U7540 ( .A(n9059), .B(g14694), .C(n12364), .Y(n9067) );
  NAND3X1 U7541 ( .A(n9057), .B(g17580), .C(n12365), .Y(n9066) );
  NAND3X1 U7542 ( .A(n9056), .B(g17711), .C(n12363), .Y(n9065) );
  OAI21X1 U7543 ( .A0(n9068), .A1(n7230), .B0(n9069), .Y(n6761) );
  AOI21X1 U7544 ( .A0(n12238), .A1(n9070), .B0(n9071), .Y(n9069) );
  AOI21X1 U7545 ( .A0(n7921), .A1(n9072), .B0(n12239), .Y(n9071) );
  NAND3X1 U7546 ( .A(n7710), .B(n7854), .C(n9073), .Y(n9072) );
  NAND2X1 U7547 ( .A(n7854), .B(n9074), .Y(n9070) );
  NAND3X1 U7548 ( .A(n9073), .B(g35), .C(n12239), .Y(n9074) );
  OAI21X1 U7549 ( .A0(n9075), .A1(n7560), .B0(n9076), .Y(n6760) );
  MX2X1 U7550 ( .A(n9077), .B(n7230), .S0(n7954), .Y(n9076) );
  NAND2X1 U7551 ( .A(n8543), .B(n7560), .Y(n9077) );
  OAI21X1 U7552 ( .A0(n12233), .A1(n9068), .B0(n9078), .Y(n6759) );
  OAI21X1 U7553 ( .A0(n9073), .A1(n8593), .B0(n12234), .Y(n9078) );
  OAI21X1 U7554 ( .A0(n12696), .A1(n9068), .B0(n9079), .Y(n6758) );
  MX2X1 U7555 ( .A(n9080), .B(n9081), .S0(n12233), .Y(n9079) );
  NAND3X1 U7556 ( .A(n7932), .B(n7560), .C(n9073), .Y(n9081) );
  AOI21X1 U7557 ( .A0(n12234), .A1(n9073), .B0(n8593), .Y(n9080) );
  OAI21X1 U7558 ( .A0(n9068), .A1(n7561), .B0(n9082), .Y(n6757) );
  MX2X1 U7559 ( .A(n9083), .B(n12696), .S0(n7953), .Y(n9082) );
  NAND2X1 U7560 ( .A(n9073), .B(n7561), .Y(n9083) );
  OR2X1 U7561 ( .A(n7965), .B(n9073), .Y(n9068) );
  NOR2X1 U7562 ( .A(n9029), .B(n9028), .Y(n9073) );
  NAND3X1 U7563 ( .A(g17604), .B(n7415), .C(n9056), .Y(n9029) );
  MX2X1 U7564 ( .A(n12231), .B(n12232), .S0(n9075), .Y(n6756) );
  OAI21X1 U7565 ( .A0(n9075), .A1(n7622), .B0(n9084), .Y(n6755) );
  MX2X1 U7566 ( .A(n9085), .B(n9086), .S0(n12231), .Y(n9084) );
  AOI21X1 U7567 ( .A0(n12232), .A1(n8543), .B0(n8593), .Y(n9086) );
  NAND3X1 U7568 ( .A(n7932), .B(n7561), .C(n8543), .Y(n9085) );
  INVX1 U7569 ( .A(n8492), .Y(n9075) );
  INVX1 U7570 ( .A(n9087), .Y(n6754) );
  AOI22X1 U7571 ( .A0(n12230), .A1(n9088), .B0(n12235), .B1(test_se), .Y(n9087) );
  NAND2X1 U7572 ( .A(n9089), .B(n9090), .Y(n6753) );
  MX2X1 U7573 ( .A(n9091), .B(n12230), .S0(n7953), .Y(n9089) );
  INVX1 U7574 ( .A(n9092), .Y(n6752) );
  AOI22X1 U7575 ( .A0(n9093), .A1(n7259), .B0(n7965), .B1(n7425), .Y(n9092) );
  OAI21X1 U7576 ( .A0(n12237), .A1(n9094), .B0(n9095), .Y(n6751) );
  OAI21X1 U7577 ( .A0(n12237), .A1(n7965), .B0(n12236), .Y(n9095) );
  INVX1 U7578 ( .A(n9088), .Y(n9094) );
  NAND2X1 U7579 ( .A(n9096), .B(n9097), .Y(n6750) );
  MX2X1 U7580 ( .A(n9098), .B(n12237), .S0(n7946), .Y(n9097) );
  AOI21X1 U7581 ( .A0(n9088), .A1(n12240), .B0(n9099), .Y(n9096) );
  NOR2X1 U7582 ( .A(n7965), .B(n12236), .Y(n9088) );
  NAND2X1 U7583 ( .A(n9100), .B(n9101), .Y(n6749) );
  MX2X1 U7584 ( .A(n9102), .B(n8534), .S0(n9103), .Y(n9101) );
  NOR2X1 U7585 ( .A(n7259), .B(n9098), .Y(n9103) );
  NAND2X1 U7586 ( .A(n12368), .B(n7932), .Y(n9102) );
  AOI22X1 U7587 ( .A0(n12358), .A1(n7905), .B0(n12362), .B1(test_se), .Y(n9100) );
  NAND2X1 U7588 ( .A(n9104), .B(n9105), .Y(n6748) );
  MX2X1 U7589 ( .A(n9106), .B(n8534), .S0(n9107), .Y(n9105) );
  NOR2X1 U7590 ( .A(n9108), .B(n9090), .Y(n9107) );
  NAND2X1 U7591 ( .A(n12355), .B(n7934), .Y(n9106) );
  AOI22X1 U7592 ( .A0(n12352), .A1(n7905), .B0(n12368), .B1(test_se), .Y(n9104) );
  NAND2X1 U7593 ( .A(n9109), .B(n9110), .Y(n6747) );
  MX2X1 U7594 ( .A(n9111), .B(n8534), .S0(n9112), .Y(n9110) );
  NOR2X1 U7595 ( .A(n9091), .B(n9108), .Y(n9112) );
  NAND2X1 U7596 ( .A(n12354), .B(n7934), .Y(n9111) );
  AOI22X1 U7597 ( .A0(n12355), .A1(n7905), .B0(n12359), .B1(test_se), .Y(n9109) );
  NAND2X1 U7598 ( .A(n9113), .B(n9114), .Y(n6746) );
  MX2X1 U7599 ( .A(n9115), .B(n8534), .S0(n9116), .Y(n9114) );
  NOR2X1 U7600 ( .A(n9117), .B(n9108), .Y(n9116) );
  NAND2X1 U7601 ( .A(n7934), .B(n7226), .Y(n9115) );
  AOI22X1 U7602 ( .A0(n12354), .A1(n7905), .B0(n12361), .B1(test_se), .Y(n9113) );
  NAND2X1 U7603 ( .A(n9118), .B(n9119), .Y(n6745) );
  AOI22X1 U7604 ( .A0(n9120), .A1(n12365), .B0(n9121), .B1(n9093), .Y(n9119)
         );
  AOI21X1 U7605 ( .A0(n9122), .A1(n9093), .B0(n7965), .Y(n9120) );
  AOI22X1 U7606 ( .A0(n12363), .A1(n7905), .B0(test_se), .B1(n7226), .Y(n9118)
         );
  NAND2X1 U7607 ( .A(n9123), .B(n9124), .Y(n6744) );
  MX2X1 U7608 ( .A(n9125), .B(n8534), .S0(n9126), .Y(n9124) );
  NOR2X1 U7609 ( .A(n9117), .B(n9098), .Y(n9126) );
  NAND2X1 U7610 ( .A(n12358), .B(n7934), .Y(n9125) );
  AOI22X1 U7611 ( .A0(n12369), .A1(n7905), .B0(n12365), .B1(test_se), .Y(n9123) );
  NAND2X1 U7612 ( .A(n9127), .B(n9128), .Y(n6743) );
  MX2X1 U7613 ( .A(n9129), .B(n8534), .S0(n9130), .Y(n9128) );
  NOR2X1 U7614 ( .A(n9131), .B(n9117), .Y(n9130) );
  INVX1 U7615 ( .A(n9093), .Y(n9117) );
  NOR2X1 U7616 ( .A(n12230), .B(n12229), .Y(n9093) );
  NAND2X1 U7617 ( .A(n12360), .B(n7934), .Y(n9129) );
  AOI22X1 U7618 ( .A0(n12361), .A1(n7905), .B0(n12358), .B1(test_se), .Y(n9127) );
  OAI21X1 U7619 ( .A0(n7934), .A1(n7790), .B0(n9132), .Y(n6742) );
  AOI22X1 U7620 ( .A0(n8492), .A1(n12371), .B0(n8893), .B1(n8543), .Y(n9132)
         );
  NOR2X1 U7621 ( .A(n7965), .B(n8543), .Y(n8492) );
  NOR2X1 U7622 ( .A(n7259), .B(n9131), .Y(n8543) );
  MX2X1 U7623 ( .A(n12371), .B(g17711), .S0(n7850), .Y(n6741) );
  INVX1 U7624 ( .A(n9133), .Y(n6740) );
  MX2X1 U7625 ( .A(n9134), .B(n7854), .S0(g13049), .Y(n9133) );
  NAND4X1 U7626 ( .A(n7817), .B(n5778), .C(n9135), .D(n7934), .Y(n9134) );
  MX2X1 U7627 ( .A(n5779), .B(g12300), .S0(g14694), .Y(n9135) );
  MX2X1 U7628 ( .A(g17604), .B(g12300), .S0(n7850), .Y(n6739) );
  MX2X1 U7629 ( .A(g12300), .B(g14694), .S0(n7851), .Y(n6738) );
  OAI21X1 U7630 ( .A0(n9136), .A1(n9137), .B0(n9138), .Y(n6736) );
  MX2X1 U7631 ( .A(n9139), .B(n7791), .S0(n7951), .Y(n9138) );
  NAND2X1 U7632 ( .A(n9136), .B(n12356), .Y(n9139) );
  INVX1 U7633 ( .A(n9140), .Y(n9136) );
  NOR2X1 U7634 ( .A(n9141), .B(n9142), .Y(n6735) );
  MX2X1 U7635 ( .A(n12380), .B(n12356), .S0(n7946), .Y(n9142) );
  NOR2X1 U7636 ( .A(n9141), .B(n7658), .Y(n6734) );
  NOR2X1 U7637 ( .A(n9137), .B(n9140), .Y(n9141) );
  NAND4X1 U7638 ( .A(g14694), .B(g17580), .C(g17711), .D(g12300), .Y(n9140) );
  INVX1 U7639 ( .A(n9143), .Y(n9137) );
  OAI21X1 U7640 ( .A0(n12382), .A1(n9144), .B0(n9145), .Y(n6733) );
  MX2X1 U7641 ( .A(n9146), .B(n7627), .S0(n7951), .Y(n9145) );
  NAND2X1 U7642 ( .A(n8357), .B(n12382), .Y(n9146) );
  INVX1 U7643 ( .A(n8358), .Y(n9144) );
  NAND2X1 U7644 ( .A(n9147), .B(n9148), .Y(n6732) );
  AOI22X1 U7645 ( .A0(n8358), .A1(n12381), .B0(n9059), .B1(n7934), .Y(n9148)
         );
  NOR2X1 U7646 ( .A(n7965), .B(n8357), .Y(n8358) );
  AOI21X1 U7647 ( .A0(n7905), .A1(n7295), .B0(n9149), .Y(n9147) );
  MX2X1 U7648 ( .A(g14694), .B(n9150), .S0(n7851), .Y(n9149) );
  NOR2X1 U7649 ( .A(n9041), .B(n9028), .Y(n9150) );
  INVX1 U7650 ( .A(n9046), .Y(n9041) );
  MX2X1 U7651 ( .A(n12381), .B(g17604), .S0(n7851), .Y(n6731) );
  NAND2X1 U7652 ( .A(n9151), .B(n9152), .Y(n6730) );
  AOI22X1 U7653 ( .A0(n8261), .A1(n9153), .B0(n9154), .B1(n7504), .Y(n9152) );
  AOI22X1 U7654 ( .A0(n12350), .A1(n7905), .B0(n12394), .B1(test_se), .Y(n9151) );
  INVX1 U7655 ( .A(n9155), .Y(n6729) );
  AOI22X1 U7656 ( .A0(n9156), .A1(n9157), .B0(n12396), .B1(test_se), .Y(n9155)
         );
  INVX1 U7657 ( .A(n8604), .Y(n9157) );
  NAND3X1 U7658 ( .A(n12549), .B(n12603), .C(n12392), .Y(n8604) );
  OAI21X1 U7659 ( .A0(n12392), .A1(n7854), .B0(n9158), .Y(n6728) );
  MX2X1 U7660 ( .A(n9159), .B(n9160), .S0(n7285), .Y(n9158) );
  NAND2X1 U7661 ( .A(n9156), .B(n12607), .Y(n9160) );
  AOI21X1 U7662 ( .A0(n7576), .A1(n7854), .B0(n7905), .Y(n9159) );
  OAI21X1 U7663 ( .A0(n7934), .A1(n7576), .B0(n9161), .Y(n6727) );
  MX2X1 U7664 ( .A(n9162), .B(n9163), .S0(n7434), .Y(n9161) );
  NAND2X1 U7665 ( .A(n9156), .B(n9162), .Y(n9163) );
  NOR2X1 U7666 ( .A(n7965), .B(n9164), .Y(n9156) );
  INVX1 U7667 ( .A(n9165), .Y(n6726) );
  AOI22X1 U7668 ( .A0(n9166), .A1(n8950), .B0(test_se), .B1(n7247), .Y(n9165)
         );
  INVX1 U7669 ( .A(n8956), .Y(n8950) );
  XOR2X1 U7670 ( .A(n9164), .B(n7250), .Y(n9166) );
  OAI21X1 U7671 ( .A0(n12609), .A1(n7934), .B0(n9167), .Y(n6725) );
  MX2X1 U7672 ( .A(n9168), .B(n9169), .S0(n7411), .Y(n9167) );
  OR2X1 U7673 ( .A(n8956), .B(n8954), .Y(n9169) );
  NAND2X1 U7674 ( .A(n7934), .B(n8953), .Y(n8956) );
  NAND2X1 U7675 ( .A(n8954), .B(n8953), .Y(n9168) );
  NAND2X1 U7676 ( .A(n8954), .B(n7363), .Y(n8953) );
  NOR2X1 U7677 ( .A(n9170), .B(n12609), .Y(n8954) );
  INVX1 U7678 ( .A(n9164), .Y(n9170) );
  NOR2X1 U7679 ( .A(n9171), .B(n7541), .Y(n9164) );
  MX2X1 U7680 ( .A(n9172), .B(n7434), .S0(n7951), .Y(n6724) );
  MX2X1 U7681 ( .A(n9171), .B(n9173), .S0(n7654), .Y(n9172) );
  NOR2X1 U7682 ( .A(n12606), .B(n9171), .Y(n9173) );
  OAI21X1 U7683 ( .A0(n9174), .A1(n7654), .B0(n9175), .Y(n6723) );
  NAND3X1 U7684 ( .A(n7934), .B(n9171), .C(n12606), .Y(n9175) );
  INVX1 U7685 ( .A(n9176), .Y(n9171) );
  AOI21X1 U7686 ( .A0(n9176), .A1(n7541), .B0(n8593), .Y(n9174) );
  NOR2X1 U7687 ( .A(n9162), .B(n12605), .Y(n9176) );
  NAND2X1 U7688 ( .A(n12607), .B(n12524), .Y(n9162) );
  MX2X1 U7689 ( .A(n12606), .B(n7431), .S0(n7851), .Y(n6722) );
  OAI21X1 U7690 ( .A0(n7934), .A1(n7624), .B0(n9177), .Y(n6721) );
  MX2X1 U7691 ( .A(n8944), .B(n8897), .S0(n7242), .Y(n9177) );
  NAND2X1 U7692 ( .A(n9178), .B(n7934), .Y(n8897) );
  INVX1 U7693 ( .A(n8896), .Y(n8944) );
  NOR2X1 U7694 ( .A(n7965), .B(n9178), .Y(n8896) );
  OAI21X1 U7695 ( .A0(n5826), .A1(n8104), .B0(n9179), .Y(n6720) );
  AOI22X1 U7696 ( .A0(n7934), .A1(n9180), .B0(n12632), .B1(n7904), .Y(n9179)
         );
  XOR2X1 U7697 ( .A(n7361), .B(n9181), .Y(n9180) );
  NAND2X1 U7698 ( .A(n9178), .B(n12632), .Y(n9181) );
  INVX1 U7699 ( .A(n8826), .Y(n9178) );
  NAND2X1 U7700 ( .A(n4770), .B(n9182), .Y(n8826) );
  NAND3X1 U7701 ( .A(n8579), .B(n7499), .C(n9183), .Y(n9182) );
  NOR2X1 U7702 ( .A(n7379), .B(n12612), .Y(n8579) );
  MX2X1 U7703 ( .A(n12633), .B(g16624), .S0(n7849), .Y(n6719) );
  INVX1 U7704 ( .A(n9184), .Y(n6718) );
  MX2X1 U7705 ( .A(n9185), .B(n7870), .S0(g14421), .Y(n9184) );
  NAND4X1 U7706 ( .A(n7837), .B(n5825), .C(n9186), .D(n7934), .Y(n9185) );
  MX2X1 U7707 ( .A(n5824), .B(g11349), .S0(g13895), .Y(n9186) );
  MX2X1 U7708 ( .A(g11349), .B(g13895), .S0(n7851), .Y(n6717) );
  MX2X1 U7709 ( .A(n12614), .B(g16718), .S0(n7851), .Y(n6716) );
  MX2X1 U7710 ( .A(g16624), .B(g11349), .S0(n7851), .Y(n6715) );
  OAI21X1 U7711 ( .A0(n524), .A1(n7870), .B0(n9187), .Y(n6713) );
  AOI21X1 U7712 ( .A0(n12584), .A1(n7904), .B0(n9188), .Y(n9187) );
  NAND2X1 U7713 ( .A(n9189), .B(n9190), .Y(n6712) );
  AOI22X1 U7714 ( .A0(n12572), .A1(n8363), .B0(n12548), .B1(n7904), .Y(n9190)
         );
  AOI21X1 U7715 ( .A0(n12583), .A1(test_se), .B0(n9191), .Y(n9189) );
  MX2X1 U7716 ( .A(n9192), .B(n9193), .S0(n9194), .Y(n9191) );
  NOR2X1 U7717 ( .A(n9195), .B(n7526), .Y(n9194) );
  NOR2X1 U7718 ( .A(n8362), .B(n7965), .Y(n9193) );
  AND2X1 U7719 ( .A(n8362), .B(n8199), .Y(n9192) );
  MX2X1 U7720 ( .A(n9196), .B(n9197), .S0(n7374), .Y(n8362) );
  NAND4X1 U7721 ( .A(n9198), .B(n9199), .C(n9200), .D(n9201), .Y(n9197) );
  OR2X1 U7722 ( .A(n9202), .B(n8205), .Y(n9201) );
  AOI22X1 U7723 ( .A0(n12565), .A1(g14451), .B0(n12567), .B1(n12566), .Y(n9202) );
  AOI22X1 U7724 ( .A0(n9203), .A1(n12569), .B0(n9204), .B1(n12568), .Y(n9200)
         );
  NOR2X1 U7725 ( .A(n5250), .B(n8208), .Y(n9204) );
  NOR2X1 U7726 ( .A(n5249), .B(n8206), .Y(n9203) );
  OR2X1 U7727 ( .A(n9205), .B(n8207), .Y(n9199) );
  AOI22X1 U7728 ( .A0(n12558), .A1(g16722), .B0(n12557), .B1(g16656), .Y(n9205) );
  MX2X1 U7729 ( .A(n9206), .B(n9207), .S0(g11388), .Y(n9198) );
  AOI21X1 U7730 ( .A0(n9208), .A1(n7386), .B0(n9209), .Y(n9207) );
  INVX1 U7731 ( .A(n9210), .Y(n9206) );
  NAND4X1 U7732 ( .A(n9211), .B(n9212), .C(n9213), .D(n9214), .Y(n9196) );
  OR2X1 U7733 ( .A(n9215), .B(n8206), .Y(n9214) );
  INVX1 U7734 ( .A(n9216), .Y(n8206) );
  AOI22X1 U7735 ( .A0(n12551), .A1(g14451), .B0(n12552), .B1(n12566), .Y(n9215) );
  AOI22X1 U7736 ( .A0(n9217), .A1(n12555), .B0(n9218), .B1(n12556), .Y(n9213)
         );
  NOR2X1 U7737 ( .A(n5250), .B(n8207), .Y(n9218) );
  NOR2X1 U7738 ( .A(n5249), .B(n8205), .Y(n9217) );
  INVX1 U7739 ( .A(n9219), .Y(n8205) );
  OR2X1 U7740 ( .A(n9220), .B(n8208), .Y(n9212) );
  INVX1 U7741 ( .A(n9208), .Y(n8208) );
  AOI22X1 U7742 ( .A0(g16722), .A1(n7279), .B0(n12554), .B1(g16656), .Y(n9220)
         );
  MX2X1 U7743 ( .A(n9221), .B(n9222), .S0(g11388), .Y(n9211) );
  AOI21X1 U7744 ( .A0(n9223), .A1(n7438), .B0(n9210), .Y(n9222) );
  NAND3X1 U7745 ( .A(n9224), .B(n9225), .C(n9226), .Y(n9210) );
  NAND3X1 U7746 ( .A(n9219), .B(g13926), .C(n12562), .Y(n9226) );
  NAND3X1 U7747 ( .A(n9216), .B(g16627), .C(n12564), .Y(n9225) );
  NAND3X1 U7748 ( .A(n9208), .B(g16744), .C(n12563), .Y(n9224) );
  INVX1 U7749 ( .A(n9209), .Y(n9221) );
  NAND3X1 U7750 ( .A(n9227), .B(n9228), .C(n9229), .Y(n9209) );
  NAND3X1 U7751 ( .A(n9223), .B(g16744), .C(n12559), .Y(n9229) );
  NAND3X1 U7752 ( .A(n9216), .B(g13926), .C(n12560), .Y(n9228) );
  NOR2X1 U7753 ( .A(n12570), .B(n12571), .Y(n9216) );
  NAND3X1 U7754 ( .A(n9219), .B(g16627), .C(n12561), .Y(n9227) );
  NAND2X1 U7755 ( .A(n9230), .B(n9231), .Y(n6711) );
  AOI22X1 U7756 ( .A0(n9232), .A1(n9233), .B0(n12673), .B1(n9234), .Y(n9231)
         );
  MX2X1 U7757 ( .A(n9235), .B(n9236), .S0(n12548), .Y(n9233) );
  NOR2X1 U7758 ( .A(n12572), .B(n9237), .Y(n9236) );
  NOR2X1 U7759 ( .A(test_se), .B(n7526), .Y(n9235) );
  NOR2X1 U7760 ( .A(n9238), .B(n9239), .Y(n9232) );
  AOI22X1 U7761 ( .A0(n12572), .A1(n7904), .B0(n12548), .B1(test_se), .Y(n9230) );
  OAI21X1 U7762 ( .A0(n9240), .A1(n7398), .B0(n9241), .Y(n6710) );
  MX2X1 U7763 ( .A(n9242), .B(n7322), .S0(n7947), .Y(n9241) );
  NAND2X1 U7764 ( .A(n8551), .B(n7398), .Y(n9242) );
  OAI21X1 U7765 ( .A0(n8721), .A1(n7398), .B0(n9243), .Y(n6709) );
  AOI21X1 U7766 ( .A0(n12544), .A1(n9234), .B0(n9244), .Y(n9243) );
  INVX1 U7767 ( .A(n9245), .Y(n9234) );
  OAI21X1 U7768 ( .A0(n9245), .A1(n7643), .B0(n9246), .Y(n6708) );
  MX2X1 U7769 ( .A(n9247), .B(n9248), .S0(n12544), .Y(n9246) );
  NOR2X1 U7770 ( .A(n9244), .B(n8593), .Y(n9248) );
  NOR3X1 U7771 ( .A(n9239), .B(n9238), .C(n7398), .Y(n9244) );
  NAND3X1 U7772 ( .A(n8199), .B(n7398), .C(n9195), .Y(n9247) );
  OAI21X1 U7773 ( .A0(n7934), .A1(n7643), .B0(n9249), .Y(n6707) );
  MX2X1 U7774 ( .A(n9245), .B(n9250), .S0(n7581), .Y(n9249) );
  NAND2X1 U7775 ( .A(n9195), .B(n8199), .Y(n9250) );
  INVX1 U7776 ( .A(n9239), .Y(n9195) );
  AOI21X1 U7777 ( .A0(n9239), .A1(n7934), .B0(n8363), .Y(n9245) );
  NAND3X1 U7778 ( .A(n9208), .B(g16656), .C(n12573), .Y(n9239) );
  NOR2X1 U7779 ( .A(n7274), .B(n7543), .Y(n9208) );
  MX2X1 U7780 ( .A(n12542), .B(n12543), .S0(n9240), .Y(n6706) );
  OAI21X1 U7781 ( .A0(n9240), .A1(n7333), .B0(n9251), .Y(n6705) );
  MX2X1 U7782 ( .A(n9252), .B(n9253), .S0(n12542), .Y(n9251) );
  AOI21X1 U7783 ( .A0(n12543), .A1(n8551), .B0(n8593), .Y(n9253) );
  NAND3X1 U7784 ( .A(n7934), .B(n7581), .C(n8551), .Y(n9252) );
  INVX1 U7785 ( .A(n8504), .Y(n9240) );
  INVX1 U7786 ( .A(n9254), .Y(n6704) );
  AOI22X1 U7787 ( .A0(n9255), .A1(n7298), .B0(n12545), .B1(test_se), .Y(n9254)
         );
  NAND2X1 U7788 ( .A(n9256), .B(n9257), .Y(n6703) );
  MX2X1 U7789 ( .A(n9258), .B(n7298), .S0(n7950), .Y(n9256) );
  INVX1 U7790 ( .A(n9259), .Y(n6702) );
  AOI22X1 U7791 ( .A0(n9260), .A1(n7220), .B0(n12534), .B1(n7965), .Y(n9259)
         );
  OAI21X1 U7792 ( .A0(n7267), .A1(n9261), .B0(n9262), .Y(n6701) );
  OAI21X1 U7793 ( .A0(n7965), .A1(n7267), .B0(n12546), .Y(n9262) );
  INVX1 U7794 ( .A(n9255), .Y(n9261) );
  NAND2X1 U7795 ( .A(n9263), .B(n9264), .Y(n6700) );
  MX2X1 U7796 ( .A(n9265), .B(n7267), .S0(n7950), .Y(n9264) );
  AOI21X1 U7797 ( .A0(n9255), .A1(n12574), .B0(n9266), .Y(n9263) );
  NOR2X1 U7798 ( .A(n7965), .B(n12546), .Y(n9255) );
  INVX1 U7799 ( .A(n9267), .Y(n6699) );
  AOI22X1 U7800 ( .A0(n12574), .A1(n7934), .B0(n12584), .B1(test_se), .Y(n9267) );
  NAND2X1 U7801 ( .A(n9268), .B(n9269), .Y(n6698) );
  MX2X1 U7802 ( .A(n9270), .B(n8534), .S0(n9271), .Y(n9269) );
  NOR2X1 U7803 ( .A(n7220), .B(n9265), .Y(n9271) );
  NAND2X1 U7804 ( .A(n12567), .B(n7934), .Y(n9270) );
  AOI22X1 U7805 ( .A0(n12558), .A1(n7904), .B0(test_se), .B1(n7386), .Y(n9268)
         );
  NAND2X1 U7806 ( .A(n9272), .B(n9273), .Y(n6697) );
  MX2X1 U7807 ( .A(n9274), .B(n8534), .S0(n9275), .Y(n9273) );
  NOR2X1 U7808 ( .A(n9276), .B(n9257), .Y(n9275) );
  NAND2X1 U7809 ( .A(n12556), .B(n7925), .Y(n9274) );
  AOI22X1 U7810 ( .A0(n12551), .A1(n7904), .B0(n12567), .B1(test_se), .Y(n9272) );
  NAND2X1 U7811 ( .A(n9277), .B(n9278), .Y(n6696) );
  MX2X1 U7812 ( .A(n9279), .B(n8534), .S0(n9280), .Y(n9278) );
  NOR2X1 U7813 ( .A(n9258), .B(n9276), .Y(n9280) );
  NAND2X1 U7814 ( .A(n12555), .B(n7923), .Y(n9279) );
  AOI22X1 U7815 ( .A0(n12556), .A1(n7904), .B0(n12560), .B1(test_se), .Y(n9277) );
  NAND2X1 U7816 ( .A(n9281), .B(n9282), .Y(n6695) );
  MX2X1 U7817 ( .A(n9283), .B(n8534), .S0(n9284), .Y(n9282) );
  NOR2X1 U7818 ( .A(n9285), .B(n9276), .Y(n9284) );
  NAND2X1 U7819 ( .A(n7923), .B(n7279), .Y(n9283) );
  AOI22X1 U7820 ( .A0(n12555), .A1(n7904), .B0(n12559), .B1(test_se), .Y(n9281) );
  NAND2X1 U7821 ( .A(n9286), .B(n9287), .Y(n6694) );
  AOI22X1 U7822 ( .A0(n9288), .A1(n12564), .B0(n9289), .B1(n9260), .Y(n9287)
         );
  AOI21X1 U7823 ( .A0(n9290), .A1(n9260), .B0(n7964), .Y(n9288) );
  AOI22X1 U7824 ( .A0(n12563), .A1(n7904), .B0(test_se), .B1(n7279), .Y(n9286)
         );
  NAND2X1 U7825 ( .A(n9291), .B(n9292), .Y(n6693) );
  MX2X1 U7826 ( .A(n9293), .B(n8534), .S0(n9294), .Y(n9292) );
  NOR2X1 U7827 ( .A(n9285), .B(n9265), .Y(n9294) );
  NAND2X1 U7828 ( .A(n12558), .B(n7923), .Y(n9293) );
  AOI22X1 U7829 ( .A0(n12569), .A1(n7904), .B0(n12564), .B1(test_se), .Y(n9291) );
  NAND2X1 U7830 ( .A(n9295), .B(n9296), .Y(n6692) );
  MX2X1 U7831 ( .A(n9297), .B(n8534), .S0(n9298), .Y(n9296) );
  NOR2X1 U7832 ( .A(n9299), .B(n9285), .Y(n9298) );
  INVX1 U7833 ( .A(n9260), .Y(n9285) );
  NOR2X1 U7834 ( .A(n7565), .B(n7298), .Y(n9260) );
  NAND2X1 U7835 ( .A(n12561), .B(n7923), .Y(n9297) );
  AOI22X1 U7836 ( .A0(n12559), .A1(n7904), .B0(n12558), .B1(test_se), .Y(n9295) );
  OAI21X1 U7837 ( .A0(n7923), .A1(n7792), .B0(n9300), .Y(n6691) );
  AOI22X1 U7838 ( .A0(n8504), .A1(n12554), .B0(n8893), .B1(n8551), .Y(n9300)
         );
  NOR2X1 U7839 ( .A(n7964), .B(n8551), .Y(n8504) );
  NOR2X1 U7840 ( .A(n7220), .B(n9299), .Y(n8551) );
  NAND2X1 U7841 ( .A(n9301), .B(n9302), .Y(n6690) );
  MX2X1 U7842 ( .A(n9303), .B(n9304), .S0(n9305), .Y(n9302) );
  INVX1 U7843 ( .A(n9188), .Y(n9304) );
  NAND2X1 U7844 ( .A(n7923), .B(n7374), .Y(n9303) );
  AOI22X1 U7845 ( .A0(n12566), .A1(n7904), .B0(n12531), .B1(test_se), .Y(n9301) );
  AOI21X1 U7846 ( .A0(n9188), .A1(n9306), .B0(n9307), .Y(n6689) );
  MX2X1 U7847 ( .A(n12530), .B(n7374), .S0(n7949), .Y(n9307) );
  NOR2X1 U7848 ( .A(n7374), .B(n7964), .Y(n9188) );
  AOI21X1 U7849 ( .A0(n9308), .A1(n9306), .B0(n12529), .Y(n6688) );
  INVX1 U7850 ( .A(n9305), .Y(n9306) );
  NAND4X1 U7851 ( .A(g16744), .B(g16627), .C(g13926), .D(g11388), .Y(n9305) );
  NOR2X1 U7852 ( .A(n7374), .B(n8593), .Y(n9308) );
  INVX1 U7853 ( .A(n9309), .Y(n6687) );
  AOI21X1 U7854 ( .A0(n7964), .A1(n12530), .B0(n9310), .Y(n9309) );
  MX2X1 U7855 ( .A(n8363), .B(n8199), .S0(n7274), .Y(n9310) );
  NOR2X1 U7856 ( .A(n9238), .B(n7964), .Y(n8199) );
  OAI21X1 U7857 ( .A0(n7984), .A1(n7870), .B0(n9311), .Y(n6686) );
  AOI21X1 U7858 ( .A0(n12528), .A1(n7903), .B0(n9312), .Y(n9311) );
  OAI21X1 U7859 ( .A0(n7870), .A1(n7748), .B0(n9313), .Y(n6685) );
  AOI22X1 U7860 ( .A0(n7923), .A1(n9314), .B0(n12500), .B1(n7903), .Y(n9313)
         );
  OAI21X1 U7861 ( .A0(n9315), .A1(n9316), .B0(n9317), .Y(n9314) );
  MX2X1 U7862 ( .A(n9318), .B(n7513), .S0(n9319), .Y(n9317) );
  NAND2X1 U7863 ( .A(n9315), .B(n9316), .Y(n9318) );
  NAND2X1 U7864 ( .A(n12501), .B(n9320), .Y(n9316) );
  NAND3X1 U7865 ( .A(n9321), .B(g16693), .C(n12525), .Y(n9320) );
  OAI21X1 U7866 ( .A0(n9322), .A1(n7620), .B0(n9323), .Y(n6684) );
  AOI21X1 U7867 ( .A0(n12500), .A1(n9324), .B0(n9325), .Y(n9323) );
  AOI21X1 U7868 ( .A0(n7921), .A1(n9326), .B0(n7513), .Y(n9325) );
  NAND3X1 U7869 ( .A(n7711), .B(n7870), .C(n9327), .Y(n9326) );
  NAND2X1 U7870 ( .A(n7870), .B(n9328), .Y(n9324) );
  NAND3X1 U7871 ( .A(g35), .B(n7513), .C(n9327), .Y(n9328) );
  OAI21X1 U7872 ( .A0(n9329), .A1(n7562), .B0(n9330), .Y(n6683) );
  MX2X1 U7873 ( .A(n9331), .B(n7620), .S0(n7949), .Y(n9330) );
  NAND2X1 U7874 ( .A(n8548), .B(n7562), .Y(n9331) );
  OAI21X1 U7875 ( .A0(n9322), .A1(n7655), .B0(n9332), .Y(n6682) );
  OAI21X1 U7876 ( .A0(n9327), .A1(n8593), .B0(n12496), .Y(n9332) );
  OAI21X1 U7877 ( .A0(n9322), .A1(n7645), .B0(n9333), .Y(n6681) );
  MX2X1 U7878 ( .A(n9334), .B(n9335), .S0(n7655), .Y(n9333) );
  NAND3X1 U7879 ( .A(n7923), .B(n7562), .C(n9327), .Y(n9335) );
  AOI21X1 U7880 ( .A0(n12496), .A1(n9327), .B0(n8593), .Y(n9334) );
  OAI21X1 U7881 ( .A0(n9322), .A1(n7563), .B0(n9336), .Y(n6680) );
  MX2X1 U7882 ( .A(n9337), .B(n7645), .S0(n7949), .Y(n9336) );
  NAND2X1 U7883 ( .A(n9327), .B(n7563), .Y(n9337) );
  INVX1 U7884 ( .A(n9338), .Y(n9327) );
  NAND2X1 U7885 ( .A(n7923), .B(n9338), .Y(n9322) );
  NAND4X1 U7886 ( .A(n12525), .B(n9321), .C(n9339), .D(g16693), .Y(n9338) );
  MX2X1 U7887 ( .A(n12494), .B(n12495), .S0(n9329), .Y(n6679) );
  OAI21X1 U7888 ( .A0(n9329), .A1(n7334), .B0(n9340), .Y(n6678) );
  MX2X1 U7889 ( .A(n9341), .B(n9342), .S0(n12494), .Y(n9340) );
  AOI21X1 U7890 ( .A0(n12495), .A1(n8548), .B0(n8593), .Y(n9342) );
  NAND3X1 U7891 ( .A(n7923), .B(n7563), .C(n8548), .Y(n9341) );
  INVX1 U7892 ( .A(n8500), .Y(n9329) );
  INVX1 U7893 ( .A(n9343), .Y(n6677) );
  AOI22X1 U7894 ( .A0(n9344), .A1(n7299), .B0(n12497), .B1(test_se), .Y(n9343)
         );
  NAND2X1 U7895 ( .A(n9345), .B(n9346), .Y(n6676) );
  MX2X1 U7896 ( .A(n9347), .B(n7299), .S0(n7948), .Y(n9345) );
  INVX1 U7897 ( .A(n9348), .Y(n6675) );
  AOI22X1 U7898 ( .A0(n9349), .A1(n7221), .B0(n12492), .B1(n7964), .Y(n9348)
         );
  OAI21X1 U7899 ( .A0(n7268), .A1(n9350), .B0(n9351), .Y(n6674) );
  OAI21X1 U7900 ( .A0(n7964), .A1(n7268), .B0(n12498), .Y(n9351) );
  INVX1 U7901 ( .A(n9344), .Y(n9350) );
  NAND2X1 U7902 ( .A(n9352), .B(n9353), .Y(n6673) );
  MX2X1 U7903 ( .A(n9354), .B(n7268), .S0(n7947), .Y(n9353) );
  AOI21X1 U7904 ( .A0(n9344), .A1(n12526), .B0(n9355), .Y(n9352) );
  NOR2X1 U7905 ( .A(n7964), .B(n12498), .Y(n9344) );
  INVX1 U7906 ( .A(n9356), .Y(n6672) );
  AOI22X1 U7907 ( .A0(n12526), .A1(n7924), .B0(n12528), .B1(test_se), .Y(n9356) );
  NAND2X1 U7908 ( .A(n9357), .B(n9358), .Y(n6671) );
  MX2X1 U7909 ( .A(n9359), .B(n8534), .S0(n9360), .Y(n9358) );
  NOR2X1 U7910 ( .A(n7221), .B(n9354), .Y(n9360) );
  NAND2X1 U7911 ( .A(n12518), .B(n7923), .Y(n9359) );
  AOI22X1 U7912 ( .A0(n12509), .A1(n7903), .B0(test_se), .B1(n7387), .Y(n9357)
         );
  NAND2X1 U7913 ( .A(n9361), .B(n9362), .Y(n6670) );
  MX2X1 U7914 ( .A(n9363), .B(n8534), .S0(n9364), .Y(n9362) );
  NOR2X1 U7915 ( .A(n9365), .B(n9346), .Y(n9364) );
  NAND2X1 U7916 ( .A(n12507), .B(n7924), .Y(n9363) );
  AOI22X1 U7917 ( .A0(n12502), .A1(n7903), .B0(n12518), .B1(test_se), .Y(n9361) );
  NAND2X1 U7918 ( .A(n9366), .B(n9367), .Y(n6669) );
  MX2X1 U7919 ( .A(n9368), .B(n8534), .S0(n9369), .Y(n9367) );
  NOR2X1 U7920 ( .A(n9347), .B(n9365), .Y(n9369) );
  NAND2X1 U7921 ( .A(n12506), .B(n7923), .Y(n9368) );
  AOI22X1 U7922 ( .A0(n12507), .A1(n7903), .B0(n12511), .B1(test_se), .Y(n9366) );
  NAND2X1 U7923 ( .A(n9370), .B(n9371), .Y(n6668) );
  MX2X1 U7924 ( .A(n9372), .B(n8534), .S0(n9373), .Y(n9371) );
  NOR2X1 U7925 ( .A(n9374), .B(n9365), .Y(n9373) );
  NAND2X1 U7926 ( .A(n7924), .B(n7280), .Y(n9372) );
  AOI22X1 U7927 ( .A0(n12506), .A1(n7903), .B0(n12510), .B1(test_se), .Y(n9370) );
  NAND2X1 U7928 ( .A(n9375), .B(n9376), .Y(n6667) );
  AOI22X1 U7929 ( .A0(n9377), .A1(n12515), .B0(n9378), .B1(n9349), .Y(n9376)
         );
  AOI21X1 U7930 ( .A0(n9379), .A1(n9349), .B0(n7964), .Y(n9377) );
  AOI22X1 U7931 ( .A0(n12514), .A1(n7903), .B0(test_se), .B1(n7280), .Y(n9375)
         );
  NAND2X1 U7932 ( .A(n9380), .B(n9381), .Y(n6666) );
  MX2X1 U7933 ( .A(n9382), .B(n8534), .S0(n9383), .Y(n9381) );
  NOR2X1 U7934 ( .A(n9374), .B(n9354), .Y(n9383) );
  NAND2X1 U7935 ( .A(n12509), .B(n7923), .Y(n9382) );
  AOI22X1 U7936 ( .A0(n12522), .A1(n7903), .B0(n12515), .B1(test_se), .Y(n9380) );
  NAND2X1 U7937 ( .A(n9384), .B(n9385), .Y(n6665) );
  MX2X1 U7938 ( .A(n9386), .B(n8534), .S0(n9387), .Y(n9385) );
  NOR2X1 U7939 ( .A(n9388), .B(n9374), .Y(n9387) );
  INVX1 U7940 ( .A(n9349), .Y(n9374) );
  NOR2X1 U7941 ( .A(n7566), .B(n7299), .Y(n9349) );
  NAND2X1 U7942 ( .A(n12512), .B(n7924), .Y(n9386) );
  AOI22X1 U7943 ( .A0(n12510), .A1(n7903), .B0(n12509), .B1(test_se), .Y(n9384) );
  OAI21X1 U7944 ( .A0(n7923), .A1(n7793), .B0(n9389), .Y(n6664) );
  AOI22X1 U7945 ( .A0(n12505), .A1(n8500), .B0(n8893), .B1(n8548), .Y(n9389)
         );
  NOR2X1 U7946 ( .A(n7964), .B(n8548), .Y(n8500) );
  NOR2X1 U7947 ( .A(n7221), .B(n9388), .Y(n8548) );
  NAND2X1 U7948 ( .A(n9390), .B(n9391), .Y(n6663) );
  AOI22X1 U7949 ( .A0(n9315), .A1(n8517), .B0(n12486), .B1(n8520), .Y(n9391)
         );
  MX2X1 U7950 ( .A(n9392), .B(n9393), .S0(n7369), .Y(n9315) );
  NAND4X1 U7951 ( .A(n9394), .B(n9395), .C(n9396), .D(n9397), .Y(n9393) );
  OR2X1 U7952 ( .A(n9398), .B(n8526), .Y(n9397) );
  AOI22X1 U7953 ( .A0(n12516), .A1(g14518), .B0(n12518), .B1(n12517), .Y(n9398) );
  AOI22X1 U7954 ( .A0(n9399), .A1(n12519), .B0(n9400), .B1(n12522), .Y(n9396)
         );
  NOR2X1 U7955 ( .A(n5247), .B(n8527), .Y(n9400) );
  NOR2X1 U7956 ( .A(n5248), .B(n8525), .Y(n9399) );
  OR2X1 U7957 ( .A(n9401), .B(n8524), .Y(n9395) );
  AOI22X1 U7958 ( .A0(n12509), .A1(g16748), .B0(n12508), .B1(g16693), .Y(n9401) );
  MX2X1 U7959 ( .A(n9402), .B(n9403), .S0(g11418), .Y(n9394) );
  AOI21X1 U7960 ( .A0(n9321), .A1(n7387), .B0(n9404), .Y(n9403) );
  INVX1 U7961 ( .A(n9405), .Y(n9402) );
  NAND4X1 U7962 ( .A(n9406), .B(n9407), .C(n9408), .D(n9409), .Y(n9392) );
  OR2X1 U7963 ( .A(n9410), .B(n8525), .Y(n9409) );
  AOI22X1 U7964 ( .A0(g16748), .A1(n7280), .B0(n12505), .B1(g16693), .Y(n9410)
         );
  AOI22X1 U7965 ( .A0(n9411), .A1(n12506), .B0(n9412), .B1(n12507), .Y(n9408)
         );
  NOR2X1 U7966 ( .A(n5248), .B(n8524), .Y(n9412) );
  NOR2X1 U7967 ( .A(n5247), .B(n8526), .Y(n9411) );
  INVX1 U7968 ( .A(n9413), .Y(n8526) );
  OR2X1 U7969 ( .A(n9414), .B(n8527), .Y(n9407) );
  INVX1 U7970 ( .A(n9415), .Y(n8527) );
  AOI22X1 U7971 ( .A0(n12502), .A1(g14518), .B0(n12503), .B1(n12517), .Y(n9414) );
  MX2X1 U7972 ( .A(n9416), .B(n9417), .S0(g11418), .Y(n9406) );
  AOI21X1 U7973 ( .A0(n9418), .A1(n7439), .B0(n9405), .Y(n9417) );
  NAND3X1 U7974 ( .A(n9419), .B(n9420), .C(n9421), .Y(n9405) );
  NAND3X1 U7975 ( .A(n9413), .B(g13966), .C(n12513), .Y(n9421) );
  NAND3X1 U7976 ( .A(n9321), .B(g16775), .C(n12514), .Y(n9420) );
  INVX1 U7977 ( .A(n8525), .Y(n9321) );
  NAND2X1 U7978 ( .A(n12520), .B(n12521), .Y(n8525) );
  NAND3X1 U7979 ( .A(n9415), .B(g16659), .C(n12515), .Y(n9419) );
  INVX1 U7980 ( .A(n9404), .Y(n9416) );
  NAND3X1 U7981 ( .A(n9422), .B(n9423), .C(n9424), .Y(n9404) );
  NAND3X1 U7982 ( .A(n9418), .B(g16775), .C(n12510), .Y(n9424) );
  INVX1 U7983 ( .A(n8524), .Y(n9418) );
  NAND3X1 U7984 ( .A(n9415), .B(g13966), .C(n12511), .Y(n9423) );
  NOR2X1 U7985 ( .A(n12520), .B(n12521), .Y(n9415) );
  NAND3X1 U7986 ( .A(n9413), .B(g16659), .C(n12512), .Y(n9422) );
  AOI22X1 U7987 ( .A0(n12505), .A1(n7903), .B0(n12517), .B1(test_se), .Y(n9390) );
  NAND2X1 U7988 ( .A(n9425), .B(n9426), .Y(n6662) );
  MX2X1 U7989 ( .A(n9427), .B(n9428), .S0(n9429), .Y(n9426) );
  INVX1 U7990 ( .A(n9312), .Y(n9428) );
  NAND2X1 U7991 ( .A(n7924), .B(n7369), .Y(n9427) );
  AOI22X1 U7992 ( .A0(n12517), .A1(n7903), .B0(n12486), .B1(test_se), .Y(n9425) );
  AOI21X1 U7993 ( .A0(n9312), .A1(n9430), .B0(n9431), .Y(n6661) );
  MX2X1 U7994 ( .A(n12485), .B(n7369), .S0(n7952), .Y(n9431) );
  NOR2X1 U7995 ( .A(n7369), .B(n7964), .Y(n9312) );
  AOI21X1 U7996 ( .A0(n9432), .A1(n9430), .B0(n12484), .Y(n6660) );
  INVX1 U7997 ( .A(n9429), .Y(n9430) );
  NAND4X1 U7998 ( .A(g16775), .B(g16659), .C(g13966), .D(g11418), .Y(n9429) );
  NOR2X1 U7999 ( .A(n8593), .B(n7369), .Y(n9432) );
  INVX1 U8000 ( .A(n9433), .Y(n6659) );
  AOI21X1 U8001 ( .A0(n7964), .A1(n12485), .B0(n9434), .Y(n9433) );
  MX2X1 U8002 ( .A(n8517), .B(n8520), .S0(n12520), .Y(n9434) );
  NOR2X1 U8003 ( .A(n9319), .B(n7964), .Y(n8517) );
  INVX1 U8004 ( .A(n9435), .Y(n6658) );
  AOI22X1 U8005 ( .A0(n12575), .A1(n7903), .B0(n12520), .B1(test_se), .Y(n9435) );
  OAI21X1 U8006 ( .A0(n9436), .A1(n9437), .B0(n9438), .Y(n6657) );
  MX2X1 U8007 ( .A(n9439), .B(n7838), .S0(n7949), .Y(n9438) );
  NAND2X1 U8008 ( .A(n12474), .B(n9436), .Y(n9439) );
  NAND2X1 U8009 ( .A(n12582), .B(n9440), .Y(n9436) );
  INVX1 U8010 ( .A(n9441), .Y(n6656) );
  AOI22X1 U8011 ( .A0(n12582), .A1(n7902), .B0(n12474), .B1(test_se), .Y(n9441) );
  NAND2X1 U8012 ( .A(n9442), .B(n7963), .Y(n6655) );
  MX2X1 U8013 ( .A(n7330), .B(n7676), .S0(n7851), .Y(n9442) );
  INVX1 U8014 ( .A(n9443), .Y(n6654) );
  AOI22X1 U8015 ( .A0(n12581), .A1(n7902), .B0(n12576), .B1(test_se), .Y(n9443) );
  AND2X1 U8016 ( .A(n8593), .B(n12578), .Y(n6653) );
  NAND2X1 U8017 ( .A(n7236), .B(n7963), .Y(n6652) );
  OAI21X1 U8018 ( .A0(n7870), .A1(n7269), .B0(n9444), .Y(n6651) );
  OAI21X1 U8019 ( .A0(n9445), .A1(n9446), .B0(n7923), .Y(n9444) );
  NAND3X1 U8020 ( .A(n12578), .B(n12581), .C(n12579), .Y(n9446) );
  NAND3X1 U8021 ( .A(n7384), .B(n7269), .C(n9447), .Y(n9445) );
  NAND2X1 U8022 ( .A(n9448), .B(n7963), .Y(n6650) );
  MX2X1 U8023 ( .A(n7384), .B(n7231), .S0(n7850), .Y(n9448) );
  NAND2X1 U8024 ( .A(n9449), .B(n7963), .Y(n6649) );
  MX2X1 U8025 ( .A(n7231), .B(n7340), .S0(n7850), .Y(n9449) );
  OR2X1 U8026 ( .A(n9450), .B(n7924), .Y(n6648) );
  MX2X1 U8027 ( .A(n12579), .B(n12483), .S0(n7850), .Y(n9450) );
  OR2X1 U8028 ( .A(n9451), .B(n7924), .Y(n6647) );
  MX2X1 U8029 ( .A(n12482), .B(n12579), .S0(n7850), .Y(n9451) );
  INVX1 U8030 ( .A(n9452), .Y(n6646) );
  AOI22X1 U8031 ( .A0(n12482), .A1(n7902), .B0(n12577), .B1(test_se), .Y(n9452) );
  OAI21X1 U8032 ( .A0(n7870), .A1(n7839), .B0(n9453), .Y(n6645) );
  AOI22X1 U8033 ( .A0(n9454), .A1(n7924), .B0(n12481), .B1(n9455), .Y(n9453)
         );
  OAI21X1 U8034 ( .A0(test_se), .A1(n9456), .B0(n7919), .Y(n9455) );
  AND2X1 U8035 ( .A(n7506), .B(n9456), .Y(n9454) );
  NAND3X1 U8036 ( .A(n7384), .B(n7269), .C(n9457), .Y(n9456) );
  OAI21X1 U8037 ( .A0(n9437), .A1(n9458), .B0(n9459), .Y(n6644) );
  MX2X1 U8038 ( .A(n9460), .B(n12580), .S0(n7947), .Y(n9459) );
  NAND2X1 U8039 ( .A(n12480), .B(n9458), .Y(n9460) );
  NAND2X1 U8040 ( .A(n9440), .B(n7384), .Y(n9458) );
  NOR2X1 U8041 ( .A(n9461), .B(n7269), .Y(n9440) );
  OAI21X1 U8042 ( .A0(n9437), .A1(n9462), .B0(n9463), .Y(n6643) );
  MX2X1 U8043 ( .A(n9464), .B(n7840), .S0(n7948), .Y(n9463) );
  NAND2X1 U8044 ( .A(n12479), .B(n9462), .Y(n9464) );
  NAND3X1 U8045 ( .A(n9457), .B(n7269), .C(n12582), .Y(n9462) );
  INVX1 U8046 ( .A(n9461), .Y(n9457) );
  NAND3X1 U8047 ( .A(n9465), .B(n7330), .C(n9447), .Y(n9461) );
  INVX1 U8048 ( .A(n9466), .Y(n9447) );
  NAND3X1 U8049 ( .A(n7676), .B(n7340), .C(n7236), .Y(n9466) );
  NAND2X1 U8050 ( .A(n12481), .B(n7924), .Y(n9437) );
  OAI21X1 U8051 ( .A0(n7870), .A1(n7712), .B0(n9467), .Y(n6642) );
  AOI21X1 U8052 ( .A0(n12474), .A1(n7902), .B0(n9468), .Y(n9467) );
  AOI21X1 U8053 ( .A0(n12471), .A1(n12473), .B0(n7963), .Y(n9468) );
  INVX1 U8054 ( .A(n9469), .Y(n6641) );
  AOI22X1 U8055 ( .A0(n12649), .A1(n7902), .B0(n12471), .B1(test_se), .Y(n9469) );
  OAI21X1 U8056 ( .A0(n7870), .A1(n7819), .B0(n9470), .Y(n6640) );
  OAI21X1 U8057 ( .A0(n12649), .A1(n12470), .B0(n7922), .Y(n9470) );
  MX2X1 U8058 ( .A(n9471), .B(n12470), .S0(n7953), .Y(n6639) );
  OR2X1 U8059 ( .A(n12472), .B(n12648), .Y(n9471) );
  OAI21X1 U8060 ( .A0(n7870), .A1(n7341), .B0(n9472), .Y(n6638) );
  AOI22X1 U8061 ( .A0(n12472), .A1(n7902), .B0(n12473), .B1(n7924), .Y(n9472)
         );
  MX2X1 U8062 ( .A(n12472), .B(g8789), .S0(n7850), .Y(n6637) );
  INVX1 U8063 ( .A(n9473), .Y(n6636) );
  MX2X1 U8064 ( .A(n7862), .B(n7826), .S0(n7850), .Y(n9473) );
  OAI21X1 U8065 ( .A0(n12468), .A1(n7870), .B0(n9474), .Y(n6635) );
  AOI22X1 U8066 ( .A0(n12467), .A1(n7902), .B0(n7924), .B1(n7749), .Y(n9474)
         );
  OAI21X1 U8067 ( .A0(n7870), .A1(n7749), .B0(n9475), .Y(n6634) );
  AOI22X1 U8068 ( .A0(n9476), .A1(n7924), .B0(n7902), .B1(n7455), .Y(n9475) );
  MX2X1 U8069 ( .A(n9477), .B(n9478), .S0(n7455), .Y(n9476) );
  XOR2X1 U8070 ( .A(n603), .B(n9479), .Y(n9478) );
  XOR2X1 U8071 ( .A(n9480), .B(n9479), .Y(n9477) );
  OAI21X1 U8072 ( .A0(n9481), .A1(n9482), .B0(n603), .Y(n9480) );
  NAND3X1 U8073 ( .A(n7825), .B(n7824), .C(n7826), .Y(n9482) );
  NAND4X1 U8074 ( .A(n5217), .B(n5215), .C(n5214), .D(n5213), .Y(n9481) );
  OAI21X1 U8075 ( .A0(n7870), .A1(n7794), .B0(n9483), .Y(n6633) );
  AOI22X1 U8076 ( .A0(n12462), .A1(n7902), .B0(n12469), .B1(n7924), .Y(n9483)
         );
  MX2X1 U8077 ( .A(n9479), .B(n12594), .S0(n7950), .Y(n6632) );
  MX2X1 U8078 ( .A(n7341), .B(n7819), .S0(n12469), .Y(n9479) );
  XOR2X1 U8079 ( .A(n7625), .B(n9484), .Y(n6631) );
  NAND2X1 U8080 ( .A(n12461), .B(n7924), .Y(n9484) );
  OAI21X1 U8081 ( .A0(n12459), .A1(n9485), .B0(n9486), .Y(n6630) );
  MX2X1 U8082 ( .A(n9487), .B(n7795), .S0(n7954), .Y(n9486) );
  NAND2X1 U8083 ( .A(n12459), .B(n9485), .Y(n9487) );
  OAI21X1 U8084 ( .A0(n12467), .A1(n9488), .B0(n9489), .Y(n6629) );
  MX2X1 U8085 ( .A(n9490), .B(n7677), .S0(n7949), .Y(n9489) );
  NAND2X1 U8086 ( .A(n12467), .B(n9488), .Y(n9490) );
  OR2X1 U8087 ( .A(n9485), .B(n7677), .Y(n9488) );
  NAND2X1 U8088 ( .A(n12460), .B(n12461), .Y(n9485) );
  NAND2X1 U8089 ( .A(n9491), .B(n9492), .Y(n6628) );
  MX2X1 U8090 ( .A(n9493), .B(n8534), .S0(n9494), .Y(n9492) );
  NOR2X1 U8091 ( .A(n7217), .B(n8864), .Y(n9494) );
  OR2X1 U8092 ( .A(n12636), .B(n12601), .Y(n8864) );
  NAND2X1 U8093 ( .A(n12617), .B(n7924), .Y(n9493) );
  AOI22X1 U8094 ( .A0(n7902), .A1(n7225), .B0(test_se), .B1(n7278), .Y(n9491)
         );
  NAND2X1 U8095 ( .A(n9495), .B(n9496), .Y(n6627) );
  MX2X1 U8096 ( .A(n9497), .B(n8534), .S0(n9498), .Y(n9496) );
  NOR2X1 U8097 ( .A(n8882), .B(n8865), .Y(n9498) );
  NAND2X1 U8098 ( .A(n7924), .B(n7278), .Y(n9497) );
  AOI22X1 U8099 ( .A0(n12617), .A1(n7902), .B0(n12616), .B1(test_se), .Y(n9495) );
  NAND2X1 U8100 ( .A(n9499), .B(n9500), .Y(n6626) );
  MX2X1 U8101 ( .A(n8534), .B(n9501), .S0(n8857), .Y(n9500) );
  OR2X1 U8102 ( .A(n8882), .B(n7217), .Y(n8857) );
  NAND2X1 U8103 ( .A(n12619), .B(n7924), .Y(n9501) );
  AOI22X1 U8104 ( .A0(n12626), .A1(n7902), .B0(n12629), .B1(test_se), .Y(n9499) );
  NAND2X1 U8105 ( .A(n9502), .B(n9503), .Y(n6625) );
  MX2X1 U8106 ( .A(n9504), .B(n8534), .S0(n9505), .Y(n9503) );
  NOR2X1 U8107 ( .A(n8865), .B(n8858), .Y(n9505) );
  NAND2X1 U8108 ( .A(n12629), .B(n7924), .Y(n9504) );
  AOI22X1 U8109 ( .A0(n12619), .A1(n7901), .B0(n12617), .B1(test_se), .Y(n9502) );
  NAND2X1 U8110 ( .A(n9506), .B(n9507), .Y(n6624) );
  MX2X1 U8111 ( .A(n9508), .B(n8534), .S0(n9509), .Y(n9507) );
  NOR2X1 U8112 ( .A(n7217), .B(n8858), .Y(n9509) );
  NAND2X1 U8113 ( .A(n12631), .B(n7924), .Y(n9508) );
  AOI22X1 U8114 ( .A0(n12620), .A1(n7901), .B0(n12624), .B1(test_se), .Y(n9506) );
  NAND2X1 U8115 ( .A(n9510), .B(n9511), .Y(n6623) );
  MX2X1 U8116 ( .A(n9512), .B(n8534), .S0(n9513), .Y(n9511) );
  NOR2X1 U8117 ( .A(n8891), .B(n8865), .Y(n9513) );
  NAND3X1 U8118 ( .A(n7301), .B(n7564), .C(n7217), .Y(n8865) );
  NAND2X1 U8119 ( .A(n12624), .B(n7925), .Y(n9512) );
  AOI22X1 U8120 ( .A0(n12631), .A1(n7901), .B0(n12619), .B1(test_se), .Y(n9510) );
  NAND2X1 U8121 ( .A(n9514), .B(n9515), .Y(n6622) );
  MX2X1 U8122 ( .A(n9516), .B(n8534), .S0(n9517), .Y(n9515) );
  NOR2X1 U8123 ( .A(n8882), .B(n8852), .Y(n9517) );
  NAND2X1 U8124 ( .A(n12627), .B(n7924), .Y(n9516) );
  AOI22X1 U8125 ( .A0(n7901), .A1(n7278), .B0(n12615), .B1(test_se), .Y(n9514)
         );
  NAND2X1 U8126 ( .A(n9518), .B(n9519), .Y(n6621) );
  MX2X1 U8127 ( .A(n9520), .B(n8534), .S0(n9521), .Y(n9519) );
  NOR2X1 U8128 ( .A(n8852), .B(n8858), .Y(n9521) );
  NAND2X1 U8129 ( .A(n12618), .B(n7924), .Y(n9520) );
  AOI22X1 U8130 ( .A0(n12629), .A1(n7901), .B0(n12627), .B1(test_se), .Y(n9518) );
  NAND2X1 U8131 ( .A(n9522), .B(n9523), .Y(n6620) );
  MX2X1 U8132 ( .A(n9524), .B(n8534), .S0(n9525), .Y(n9523) );
  NOR2X1 U8133 ( .A(n8891), .B(n8852), .Y(n9525) );
  NAND2X1 U8134 ( .A(n12592), .B(n7564), .Y(n8852) );
  NAND2X1 U8135 ( .A(n12623), .B(n7924), .Y(n9524) );
  AOI22X1 U8136 ( .A0(n12624), .A1(n7901), .B0(n12618), .B1(test_se), .Y(n9522) );
  NAND2X1 U8137 ( .A(n9526), .B(n9527), .Y(n6619) );
  MX2X1 U8138 ( .A(n9528), .B(n8534), .S0(n9529), .Y(n9527) );
  NOR2X1 U8139 ( .A(n8853), .B(n8882), .Y(n9529) );
  NAND2X1 U8140 ( .A(n12601), .B(n7480), .Y(n8882) );
  NAND2X1 U8141 ( .A(n12625), .B(n7925), .Y(n9528) );
  AOI22X1 U8142 ( .A0(n12627), .A1(n7901), .B0(n12613), .B1(test_se), .Y(n9526) );
  NAND2X1 U8143 ( .A(n9530), .B(n9531), .Y(n6618) );
  MX2X1 U8144 ( .A(n9532), .B(n8534), .S0(n9533), .Y(n9531) );
  NOR2X1 U8145 ( .A(n8853), .B(n8858), .Y(n9533) );
  OR2X1 U8146 ( .A(n7480), .B(n12601), .Y(n8858) );
  NAND2X1 U8147 ( .A(n12628), .B(n7924), .Y(n9532) );
  AOI22X1 U8148 ( .A0(n12618), .A1(n7901), .B0(n12625), .B1(test_se), .Y(n9530) );
  NAND2X1 U8149 ( .A(n9534), .B(n9535), .Y(n6617) );
  MX2X1 U8150 ( .A(n9536), .B(n8534), .S0(n9537), .Y(n9535) );
  NOR2X1 U8151 ( .A(n8891), .B(n8853), .Y(n9537) );
  NAND2X1 U8152 ( .A(n12591), .B(n7301), .Y(n8853) );
  NAND2X1 U8153 ( .A(n12601), .B(n12636), .Y(n8891) );
  NAND2X1 U8154 ( .A(n12622), .B(n7925), .Y(n9536) );
  AOI22X1 U8155 ( .A0(n12623), .A1(n7901), .B0(n12628), .B1(test_se), .Y(n9534) );
  OAI21X1 U8156 ( .A0(n8534), .A1(n9538), .B0(n9539), .Y(n6616) );
  MX2X1 U8157 ( .A(n9540), .B(n7507), .S0(n7954), .Y(n9539) );
  NAND2X1 U8158 ( .A(n12551), .B(n9538), .Y(n9540) );
  OR2X1 U8159 ( .A(n9541), .B(n9276), .Y(n9538) );
  NAND2X1 U8160 ( .A(n9542), .B(n9543), .Y(n6615) );
  MX2X1 U8161 ( .A(n9544), .B(n8534), .S0(n9545), .Y(n9543) );
  NOR2X1 U8162 ( .A(n7220), .B(n9276), .Y(n9545) );
  NAND2X1 U8163 ( .A(n7507), .B(n7267), .Y(n9276) );
  NAND2X1 U8164 ( .A(n12552), .B(n7925), .Y(n9544) );
  AOI22X1 U8165 ( .A0(n7901), .A1(n7279), .B0(test_se), .B1(n7438), .Y(n9542)
         );
  NAND2X1 U8166 ( .A(n9546), .B(n9547), .Y(n6614) );
  AOI22X1 U8167 ( .A0(n9548), .A1(n7925), .B0(n9549), .B1(n9289), .Y(n9547) );
  AOI21X1 U8168 ( .A0(n9549), .A1(n9290), .B0(n12553), .Y(n9548) );
  INVX1 U8169 ( .A(n9541), .Y(n9549) );
  AOI22X1 U8170 ( .A0(n12552), .A1(n7901), .B0(n12551), .B1(test_se), .Y(n9546) );
  NAND2X1 U8171 ( .A(n9550), .B(n9551), .Y(n6613) );
  AOI22X1 U8172 ( .A0(n9552), .A1(n12557), .B0(n9289), .B1(n12546), .Y(n9551)
         );
  NOR2X1 U8173 ( .A(n9266), .B(n7962), .Y(n9552) );
  AND2X1 U8174 ( .A(n9290), .B(n12546), .Y(n9266) );
  AOI22X1 U8175 ( .A0(n12564), .A1(n7901), .B0(n12565), .B1(test_se), .Y(n9550) );
  NAND2X1 U8176 ( .A(n9553), .B(n9554), .Y(n6612) );
  MX2X1 U8177 ( .A(n9555), .B(n8534), .S0(n9556), .Y(n9554) );
  NOR2X1 U8178 ( .A(n9265), .B(n9541), .Y(n9556) );
  NAND2X1 U8179 ( .A(n12565), .B(n7925), .Y(n9555) );
  AOI22X1 U8180 ( .A0(n12557), .A1(n7900), .B0(n12552), .B1(test_se), .Y(n9553) );
  NAND2X1 U8181 ( .A(n9557), .B(n9558), .Y(n6611) );
  MX2X1 U8182 ( .A(n9559), .B(n8534), .S0(n9560), .Y(n9558) );
  NOR2X1 U8183 ( .A(n9299), .B(n9541), .Y(n9560) );
  NAND3X1 U8184 ( .A(n7298), .B(n7565), .C(n7220), .Y(n9541) );
  NAND2X1 U8185 ( .A(n7925), .B(n7386), .Y(n9559) );
  AOI22X1 U8186 ( .A0(n12567), .A1(n7900), .B0(n12557), .B1(test_se), .Y(n9557) );
  NAND2X1 U8187 ( .A(n9561), .B(n9562), .Y(n6610) );
  AOI22X1 U8188 ( .A0(n9563), .A1(n12562), .B0(n9289), .B1(n9564), .Y(n9562)
         );
  AOI21X1 U8189 ( .A0(n9564), .A1(n9290), .B0(n7962), .Y(n9563) );
  AOI22X1 U8190 ( .A0(n7900), .A1(n7438), .B0(n12556), .B1(test_se), .Y(n9561)
         );
  NAND2X1 U8191 ( .A(n9565), .B(n9566), .Y(n6609) );
  MX2X1 U8192 ( .A(n9567), .B(n8534), .S0(n9568), .Y(n9566) );
  NOR2X1 U8193 ( .A(n9265), .B(n9257), .Y(n9568) );
  NAND2X1 U8194 ( .A(n12568), .B(n7925), .Y(n9567) );
  AOI22X1 U8195 ( .A0(n12565), .A1(n7900), .B0(n12562), .B1(test_se), .Y(n9565) );
  NAND2X1 U8196 ( .A(n9569), .B(n9570), .Y(n6608) );
  MX2X1 U8197 ( .A(n9571), .B(n8534), .S0(n9572), .Y(n9570) );
  NOR2X1 U8198 ( .A(n9299), .B(n9257), .Y(n9572) );
  INVX1 U8199 ( .A(n9564), .Y(n9257) );
  NOR2X1 U8200 ( .A(n7298), .B(n12534), .Y(n9564) );
  NAND2X1 U8201 ( .A(n12560), .B(n7925), .Y(n9571) );
  AOI22X1 U8202 ( .A0(n7900), .A1(n7386), .B0(n12568), .B1(test_se), .Y(n9569)
         );
  NAND2X1 U8203 ( .A(n9573), .B(n9574), .Y(n6607) );
  AOI22X1 U8204 ( .A0(n9575), .A1(n12563), .B0(n9289), .B1(n9576), .Y(n9574)
         );
  AND2X1 U8205 ( .A(n9290), .B(n8893), .Y(n9289) );
  AOI21X1 U8206 ( .A0(n9290), .A1(n9576), .B0(n7962), .Y(n9575) );
  NOR2X1 U8207 ( .A(n7267), .B(n12574), .Y(n9290) );
  AOI22X1 U8208 ( .A0(n12562), .A1(n7900), .B0(n12555), .B1(test_se), .Y(n9573) );
  NAND2X1 U8209 ( .A(n9577), .B(n9578), .Y(n6606) );
  MX2X1 U8210 ( .A(n9579), .B(n8534), .S0(n9580), .Y(n9578) );
  NOR2X1 U8211 ( .A(n9258), .B(n9265), .Y(n9580) );
  NAND2X1 U8212 ( .A(n12574), .B(n7267), .Y(n9265) );
  NAND2X1 U8213 ( .A(n12569), .B(n7925), .Y(n9579) );
  AOI22X1 U8214 ( .A0(n12568), .A1(n7900), .B0(n12563), .B1(test_se), .Y(n9577) );
  NAND2X1 U8215 ( .A(n9581), .B(n9582), .Y(n6605) );
  MX2X1 U8216 ( .A(n9583), .B(n8534), .S0(n9584), .Y(n9582) );
  NOR2X1 U8217 ( .A(n9299), .B(n9258), .Y(n9584) );
  INVX1 U8218 ( .A(n9576), .Y(n9258) );
  NOR2X1 U8219 ( .A(n7565), .B(n12535), .Y(n9576) );
  NAND2X1 U8220 ( .A(n12547), .B(n12574), .Y(n9299) );
  NAND2X1 U8221 ( .A(n12559), .B(n7925), .Y(n9583) );
  AOI22X1 U8222 ( .A0(n12560), .A1(n7900), .B0(n12569), .B1(test_se), .Y(n9581) );
  OAI21X1 U8223 ( .A0(n8534), .A1(n9585), .B0(n9586), .Y(n6604) );
  MX2X1 U8224 ( .A(n9587), .B(n7508), .S0(n7950), .Y(n9586) );
  NAND2X1 U8225 ( .A(n12502), .B(n9585), .Y(n9587) );
  OR2X1 U8226 ( .A(n9588), .B(n9365), .Y(n9585) );
  NAND2X1 U8227 ( .A(n9589), .B(n9590), .Y(n6603) );
  MX2X1 U8228 ( .A(n9591), .B(n8534), .S0(n9592), .Y(n9590) );
  NOR2X1 U8229 ( .A(n7221), .B(n9365), .Y(n9592) );
  NAND2X1 U8230 ( .A(n7508), .B(n7268), .Y(n9365) );
  NAND2X1 U8231 ( .A(n12503), .B(n7925), .Y(n9591) );
  AOI22X1 U8232 ( .A0(n7900), .A1(n7280), .B0(test_se), .B1(n7439), .Y(n9589)
         );
  NAND2X1 U8233 ( .A(n9593), .B(n9594), .Y(n6602) );
  AOI22X1 U8234 ( .A0(n9595), .A1(n7925), .B0(n9596), .B1(n9378), .Y(n9594) );
  AOI21X1 U8235 ( .A0(n9596), .A1(n9379), .B0(n12504), .Y(n9595) );
  INVX1 U8236 ( .A(n9588), .Y(n9596) );
  AOI22X1 U8237 ( .A0(n12503), .A1(n7900), .B0(n12502), .B1(test_se), .Y(n9593) );
  NAND2X1 U8238 ( .A(n9597), .B(n9598), .Y(n6601) );
  AOI22X1 U8239 ( .A0(n9599), .A1(n12508), .B0(n9378), .B1(n12498), .Y(n9598)
         );
  NOR2X1 U8240 ( .A(n9355), .B(n7962), .Y(n9599) );
  AND2X1 U8241 ( .A(n9379), .B(n12498), .Y(n9355) );
  AOI22X1 U8242 ( .A0(n12515), .A1(n7900), .B0(n12516), .B1(test_se), .Y(n9597) );
  NAND2X1 U8243 ( .A(n9600), .B(n9601), .Y(n6600) );
  MX2X1 U8244 ( .A(n9602), .B(n8534), .S0(n9603), .Y(n9601) );
  NOR2X1 U8245 ( .A(n9354), .B(n9588), .Y(n9603) );
  NAND2X1 U8246 ( .A(n12516), .B(n7925), .Y(n9602) );
  AOI22X1 U8247 ( .A0(n12508), .A1(n7900), .B0(n12503), .B1(test_se), .Y(n9600) );
  NAND2X1 U8248 ( .A(n9604), .B(n9605), .Y(n6599) );
  MX2X1 U8249 ( .A(n9606), .B(n8534), .S0(n9607), .Y(n9605) );
  NOR2X1 U8250 ( .A(n9388), .B(n9588), .Y(n9607) );
  NAND3X1 U8251 ( .A(n7299), .B(n7566), .C(n7221), .Y(n9588) );
  NAND2X1 U8252 ( .A(n7925), .B(n7387), .Y(n9606) );
  AOI22X1 U8253 ( .A0(n12518), .A1(n7899), .B0(n12508), .B1(test_se), .Y(n9604) );
  NAND2X1 U8254 ( .A(n9608), .B(n9609), .Y(n6598) );
  AOI22X1 U8255 ( .A0(n9610), .A1(n12513), .B0(n9378), .B1(n9611), .Y(n9609)
         );
  AOI21X1 U8256 ( .A0(n9611), .A1(n9379), .B0(n7962), .Y(n9610) );
  AOI22X1 U8257 ( .A0(n7899), .A1(n7439), .B0(n12507), .B1(test_se), .Y(n9608)
         );
  NAND2X1 U8258 ( .A(n9612), .B(n9613), .Y(n6597) );
  MX2X1 U8259 ( .A(n9614), .B(n8534), .S0(n9615), .Y(n9613) );
  NOR2X1 U8260 ( .A(n9354), .B(n9346), .Y(n9615) );
  NAND2X1 U8261 ( .A(n12519), .B(n7925), .Y(n9614) );
  AOI22X1 U8262 ( .A0(n12516), .A1(n7899), .B0(n12513), .B1(test_se), .Y(n9612) );
  NAND2X1 U8263 ( .A(n9616), .B(n9617), .Y(n6596) );
  MX2X1 U8264 ( .A(n9618), .B(n8534), .S0(n9619), .Y(n9617) );
  NOR2X1 U8265 ( .A(n9388), .B(n9346), .Y(n9619) );
  INVX1 U8266 ( .A(n9611), .Y(n9346) );
  NOR2X1 U8267 ( .A(n7299), .B(n12492), .Y(n9611) );
  NAND2X1 U8268 ( .A(n12511), .B(n7925), .Y(n9618) );
  AOI22X1 U8269 ( .A0(n7899), .A1(n7387), .B0(n12519), .B1(test_se), .Y(n9616)
         );
  NAND2X1 U8270 ( .A(n9620), .B(n9621), .Y(n6595) );
  AOI22X1 U8271 ( .A0(n9622), .A1(n12514), .B0(n9378), .B1(n9623), .Y(n9621)
         );
  AND2X1 U8272 ( .A(n9379), .B(n8893), .Y(n9378) );
  AOI21X1 U8273 ( .A0(n9379), .A1(n9623), .B0(n7962), .Y(n9622) );
  NOR2X1 U8274 ( .A(n7268), .B(n12526), .Y(n9379) );
  AOI22X1 U8275 ( .A0(n12513), .A1(n7899), .B0(n12506), .B1(test_se), .Y(n9620) );
  NAND2X1 U8276 ( .A(n9624), .B(n9625), .Y(n6594) );
  MX2X1 U8277 ( .A(n9626), .B(n8534), .S0(n9627), .Y(n9625) );
  NOR2X1 U8278 ( .A(n9347), .B(n9354), .Y(n9627) );
  NAND2X1 U8279 ( .A(n12526), .B(n7268), .Y(n9354) );
  NAND2X1 U8280 ( .A(n12522), .B(n7925), .Y(n9626) );
  AOI22X1 U8281 ( .A0(n12519), .A1(n7899), .B0(n12514), .B1(test_se), .Y(n9624) );
  NAND2X1 U8282 ( .A(n9628), .B(n9629), .Y(n6593) );
  MX2X1 U8283 ( .A(n9630), .B(n8534), .S0(n9631), .Y(n9629) );
  NOR2X1 U8284 ( .A(n9388), .B(n9347), .Y(n9631) );
  INVX1 U8285 ( .A(n9623), .Y(n9347) );
  NOR2X1 U8286 ( .A(n7566), .B(n12493), .Y(n9623) );
  NAND2X1 U8287 ( .A(n12499), .B(n12526), .Y(n9388) );
  NAND2X1 U8288 ( .A(n12510), .B(n7925), .Y(n9630) );
  AOI22X1 U8289 ( .A0(n12511), .A1(n7899), .B0(n12522), .B1(test_se), .Y(n9628) );
  OAI21X1 U8290 ( .A0(n8534), .A1(n9632), .B0(n9633), .Y(n6592) );
  MX2X1 U8291 ( .A(n9634), .B(n7481), .S0(n7953), .Y(n9633) );
  NAND2X1 U8292 ( .A(n12352), .B(n9632), .Y(n9634) );
  OR2X1 U8293 ( .A(n9635), .B(n9108), .Y(n9632) );
  NAND2X1 U8294 ( .A(n9636), .B(n9637), .Y(n6591) );
  MX2X1 U8295 ( .A(n9638), .B(n8534), .S0(n9639), .Y(n9637) );
  NOR2X1 U8296 ( .A(n7259), .B(n9108), .Y(n9639) );
  NAND2X1 U8297 ( .A(n12237), .B(n7481), .Y(n9108) );
  NAND2X1 U8298 ( .A(n12353), .B(n7925), .Y(n9638) );
  AOI22X1 U8299 ( .A0(n7899), .A1(n7226), .B0(test_se), .B1(n7440), .Y(n9636)
         );
  NAND2X1 U8300 ( .A(n9640), .B(n9641), .Y(n6590) );
  AOI22X1 U8301 ( .A0(n9642), .A1(n7925), .B0(n9643), .B1(n9121), .Y(n9641) );
  AOI21X1 U8302 ( .A0(n9643), .A1(n9122), .B0(n12351), .Y(n9642) );
  INVX1 U8303 ( .A(n9635), .Y(n9643) );
  AOI22X1 U8304 ( .A0(n12353), .A1(n7899), .B0(n12352), .B1(test_se), .Y(n9640) );
  NAND2X1 U8305 ( .A(n9644), .B(n9645), .Y(n6589) );
  AOI22X1 U8306 ( .A0(n9646), .A1(n12357), .B0(n9121), .B1(n12236), .Y(n9645)
         );
  NOR2X1 U8307 ( .A(n9099), .B(n7962), .Y(n9646) );
  AND2X1 U8308 ( .A(n9122), .B(n12236), .Y(n9099) );
  AOI22X1 U8309 ( .A0(n12365), .A1(n7899), .B0(n12366), .B1(test_se), .Y(n9644) );
  NAND2X1 U8310 ( .A(n9647), .B(n9648), .Y(n6588) );
  MX2X1 U8311 ( .A(n9649), .B(n8534), .S0(n9650), .Y(n9648) );
  NOR2X1 U8312 ( .A(n9098), .B(n9635), .Y(n9650) );
  NAND2X1 U8313 ( .A(n12366), .B(n7925), .Y(n9649) );
  AOI22X1 U8314 ( .A0(n12357), .A1(n7899), .B0(n12353), .B1(test_se), .Y(n9647) );
  NAND2X1 U8315 ( .A(n9651), .B(n9652), .Y(n6587) );
  MX2X1 U8316 ( .A(n9653), .B(n8534), .S0(n9654), .Y(n9652) );
  NOR2X1 U8317 ( .A(n9131), .B(n9635), .Y(n9654) );
  NAND3X1 U8318 ( .A(n12230), .B(n7259), .C(n12229), .Y(n9635) );
  NAND2X1 U8319 ( .A(n12362), .B(n7925), .Y(n9653) );
  AOI22X1 U8320 ( .A0(n12368), .A1(n7899), .B0(n12357), .B1(test_se), .Y(n9651) );
  NAND2X1 U8321 ( .A(n9655), .B(n9656), .Y(n6586) );
  AOI22X1 U8322 ( .A0(n9657), .A1(n12364), .B0(n9121), .B1(n9658), .Y(n9656)
         );
  AOI21X1 U8323 ( .A0(n9658), .A1(n9122), .B0(n7961), .Y(n9657) );
  AOI22X1 U8324 ( .A0(n7898), .A1(n7440), .B0(n12355), .B1(test_se), .Y(n9655)
         );
  NAND2X1 U8325 ( .A(n9659), .B(n9660), .Y(n6585) );
  MX2X1 U8326 ( .A(n9661), .B(n8534), .S0(n9662), .Y(n9660) );
  NOR2X1 U8327 ( .A(n9098), .B(n9090), .Y(n9662) );
  NAND2X1 U8328 ( .A(n12370), .B(n7926), .Y(n9661) );
  AOI22X1 U8329 ( .A0(n12366), .A1(n7898), .B0(n12364), .B1(test_se), .Y(n9659) );
  NAND2X1 U8330 ( .A(n9663), .B(n9664), .Y(n6584) );
  MX2X1 U8331 ( .A(n9665), .B(n8534), .S0(n9666), .Y(n9664) );
  NOR2X1 U8332 ( .A(n9131), .B(n9090), .Y(n9666) );
  INVX1 U8333 ( .A(n9658), .Y(n9090) );
  NOR2X1 U8334 ( .A(n7425), .B(n12230), .Y(n9658) );
  NAND2X1 U8335 ( .A(n12359), .B(n7926), .Y(n9665) );
  AOI22X1 U8336 ( .A0(n12362), .A1(n7898), .B0(n12370), .B1(test_se), .Y(n9663) );
  NAND2X1 U8337 ( .A(n9667), .B(n9668), .Y(n6583) );
  AOI22X1 U8338 ( .A0(n9669), .A1(n12363), .B0(n9121), .B1(n9670), .Y(n9668)
         );
  AND2X1 U8339 ( .A(n9122), .B(n8893), .Y(n9121) );
  AOI21X1 U8340 ( .A0(n9122), .A1(n9670), .B0(n7951), .Y(n9669) );
  INVX1 U8341 ( .A(n9091), .Y(n9670) );
  NOR2X1 U8342 ( .A(n12240), .B(n12237), .Y(n9122) );
  AOI22X1 U8343 ( .A0(n12364), .A1(n7898), .B0(n12354), .B1(test_se), .Y(n9667) );
  NAND2X1 U8344 ( .A(n9671), .B(n9672), .Y(n6582) );
  MX2X1 U8345 ( .A(n9673), .B(n8534), .S0(n9674), .Y(n9672) );
  NOR2X1 U8346 ( .A(n9091), .B(n9098), .Y(n9674) );
  NAND2X1 U8347 ( .A(n12237), .B(n12240), .Y(n9098) );
  NAND2X1 U8348 ( .A(n12369), .B(n7926), .Y(n9673) );
  AOI22X1 U8349 ( .A0(n12370), .A1(n7898), .B0(n12363), .B1(test_se), .Y(n9671) );
  NAND2X1 U8350 ( .A(n9675), .B(n9676), .Y(n6581) );
  MX2X1 U8351 ( .A(n9677), .B(n8534), .S0(n9678), .Y(n9676) );
  NOR2X1 U8352 ( .A(n9131), .B(n9091), .Y(n9678) );
  NAND2X1 U8353 ( .A(n12230), .B(n7425), .Y(n9091) );
  OR2X1 U8354 ( .A(n7481), .B(n12237), .Y(n9131) );
  NAND2X1 U8355 ( .A(n12361), .B(n7926), .Y(n9677) );
  AOI22X1 U8356 ( .A0(n12359), .A1(n7898), .B0(n12369), .B1(test_se), .Y(n9675) );
  OAI21X1 U8357 ( .A0(n7870), .A1(n7539), .B0(n9679), .Y(n6580) );
  AOI22X1 U8358 ( .A0(n9680), .A1(n5677), .B0(n12466), .B1(n7898), .Y(n9679)
         );
  NOR2X1 U8359 ( .A(n12458), .B(n7960), .Y(n9680) );
  MX2X1 U8360 ( .A(n9681), .B(n12458), .S0(n7946), .Y(n6579) );
  OR2X1 U8361 ( .A(n12462), .B(n12463), .Y(n9681) );
  INVX1 U8362 ( .A(n9682), .Y(n6578) );
  AOI22X1 U8363 ( .A0(n9683), .A1(n9684), .B0(n12653), .B1(test_se), .Y(n9682)
         );
  XOR2X1 U8364 ( .A(n7375), .B(n9685), .Y(n9683) );
  OAI21X1 U8365 ( .A0(n12541), .A1(n7926), .B0(n9686), .Y(n6577) );
  MX2X1 U8366 ( .A(n9687), .B(n9688), .S0(n7252), .Y(n9686) );
  NAND2X1 U8367 ( .A(n9684), .B(n9687), .Y(n9688) );
  INVX1 U8368 ( .A(n9689), .Y(n6576) );
  AOI22X1 U8369 ( .A0(n7364), .A1(n9684), .B0(n7252), .B1(n9690), .Y(n9689) );
  OAI21X1 U8370 ( .A0(n9687), .A1(n8972), .B0(n8721), .Y(n9690) );
  NAND2X1 U8371 ( .A(n9685), .B(n7375), .Y(n9687) );
  NOR2X1 U8372 ( .A(n7959), .B(n8972), .Y(n9684) );
  INVX1 U8373 ( .A(n8988), .Y(n8972) );
  NAND3X1 U8374 ( .A(n7252), .B(n7364), .C(n9685), .Y(n8988) );
  NOR2X1 U8375 ( .A(n9691), .B(n12451), .Y(n9685) );
  OAI21X1 U8376 ( .A0(n12539), .A1(n7870), .B0(n9692), .Y(n6575) );
  AOI22X1 U8377 ( .A0(n9693), .A1(n7926), .B0(n7898), .B1(n7245), .Y(n9692) );
  XOR2X1 U8378 ( .A(n9694), .B(n12453), .Y(n9693) );
  OAI21X1 U8379 ( .A0(n7409), .A1(n9695), .B0(n9696), .Y(n6574) );
  MX2X1 U8380 ( .A(n9697), .B(n12453), .S0(n7954), .Y(n9696) );
  NAND2X1 U8381 ( .A(n9695), .B(n7409), .Y(n9697) );
  OAI21X1 U8382 ( .A0(n7353), .A1(n9691), .B0(n9698), .Y(n6573) );
  MX2X1 U8383 ( .A(n9699), .B(n12452), .S0(n7948), .Y(n9698) );
  NAND2X1 U8384 ( .A(n9691), .B(n7353), .Y(n9699) );
  OR2X1 U8385 ( .A(n9695), .B(n12452), .Y(n9691) );
  OR2X1 U8386 ( .A(n9694), .B(n12453), .Y(n9695) );
  NAND3X1 U8387 ( .A(n7413), .B(n7277), .C(n12456), .Y(n9694) );
  NAND2X1 U8388 ( .A(n9700), .B(n9701), .Y(n6572) );
  AOI22X1 U8389 ( .A0(n8520), .A1(n12521), .B0(n9413), .B1(n7926), .Y(n9701)
         );
  NOR2X1 U8390 ( .A(n7542), .B(n12520), .Y(n9413) );
  NOR2X1 U8391 ( .A(n7957), .B(n9339), .Y(n8520) );
  INVX1 U8392 ( .A(n9319), .Y(n9339) );
  AOI21X1 U8393 ( .A0(n12520), .A1(n7898), .B0(n9702), .Y(n9700) );
  MX2X1 U8394 ( .A(g13966), .B(n9703), .S0(n7850), .Y(n9702) );
  NOR2X1 U8395 ( .A(n9319), .B(n8524), .Y(n9703) );
  NAND2X1 U8396 ( .A(n12520), .B(n7542), .Y(n8524) );
  NAND2X1 U8397 ( .A(n12524), .B(n9704), .Y(n9319) );
  NAND3X1 U8398 ( .A(n12523), .B(n8340), .C(n9183), .Y(n9704) );
  NOR2X1 U8399 ( .A(n12612), .B(n12611), .Y(n8340) );
  MX2X1 U8400 ( .A(n12521), .B(g16693), .S0(n7850), .Y(n6571) );
  INVX1 U8401 ( .A(n9705), .Y(n6570) );
  MX2X1 U8402 ( .A(n9706), .B(n7870), .S0(g14518), .Y(n9705) );
  NAND4X1 U8403 ( .A(n7829), .B(n5720), .C(n9707), .D(n7926), .Y(n9706) );
  MX2X1 U8404 ( .A(n5719), .B(g11418), .S0(g13966), .Y(n9707) );
  MX2X1 U8405 ( .A(g11418), .B(g13966), .S0(n7849), .Y(n6569) );
  MX2X1 U8406 ( .A(n12505), .B(g16775), .S0(n7849), .Y(n6568) );
  MX2X1 U8407 ( .A(g16693), .B(g11418), .S0(n7851), .Y(n6567) );
  NAND2X1 U8408 ( .A(n9708), .B(n9709), .Y(n6565) );
  AOI22X1 U8409 ( .A0(n9219), .A1(n7926), .B0(n8363), .B1(n12570), .Y(n9709)
         );
  INVX1 U8410 ( .A(n8202), .Y(n8363) );
  NAND2X1 U8411 ( .A(n7926), .B(n9238), .Y(n8202) );
  NOR2X1 U8412 ( .A(n7543), .B(n12571), .Y(n9219) );
  AOI21X1 U8413 ( .A0(n12571), .A1(n7898), .B0(n9710), .Y(n9708) );
  MX2X1 U8414 ( .A(g13926), .B(n9711), .S0(n7849), .Y(n9710) );
  NOR2X1 U8415 ( .A(n9238), .B(n8207), .Y(n9711) );
  INVX1 U8416 ( .A(n9223), .Y(n8207) );
  NOR2X1 U8417 ( .A(n7274), .B(n12570), .Y(n9223) );
  NAND2X1 U8418 ( .A(n4771), .B(n9712), .Y(n9238) );
  NAND3X1 U8419 ( .A(n12550), .B(n8523), .C(n9183), .Y(n9712) );
  NOR2X1 U8420 ( .A(n7247), .B(n12611), .Y(n8523) );
  MX2X1 U8421 ( .A(n12570), .B(g16656), .S0(n7849), .Y(n6564) );
  INVX1 U8422 ( .A(n9713), .Y(n6563) );
  MX2X1 U8423 ( .A(n9714), .B(n7870), .S0(g14451), .Y(n9713) );
  NAND4X1 U8424 ( .A(n7833), .B(n5746), .C(n9715), .D(n7926), .Y(n9714) );
  MX2X1 U8425 ( .A(n5745), .B(g11388), .S0(g13926), .Y(n9715) );
  MX2X1 U8426 ( .A(g11388), .B(g13926), .S0(n7849), .Y(n6562) );
  MX2X1 U8427 ( .A(n12554), .B(g16744), .S0(n7849), .Y(n6561) );
  MX2X1 U8428 ( .A(g16656), .B(g11388), .S0(n7849), .Y(n6560) );
  NAND2X1 U8429 ( .A(n9716), .B(n9717), .Y(n6558) );
  AOI22X1 U8430 ( .A0(n9718), .A1(n7926), .B0(n7898), .B1(n7248), .Y(n9717) );
  AOI21X1 U8431 ( .A0(n8349), .A1(n12305), .B0(n9719), .Y(n9716) );
  MX2X1 U8432 ( .A(g14828), .B(n9720), .S0(n7849), .Y(n9719) );
  NOR2X1 U8433 ( .A(n9721), .B(n8255), .Y(n9720) );
  MX2X1 U8434 ( .A(n12305), .B(g17722), .S0(n7849), .Y(n6557) );
  INVX1 U8435 ( .A(n9722), .Y(n6556) );
  MX2X1 U8436 ( .A(n9723), .B(n7870), .S0(g13099), .Y(n9722) );
  NAND4X1 U8437 ( .A(n7805), .B(n5672), .C(n9724), .D(n7926), .Y(n9723) );
  MX2X1 U8438 ( .A(n5671), .B(g12470), .S0(g14828), .Y(n9724) );
  NAND2X1 U8439 ( .A(n9725), .B(n9726), .Y(n6555) );
  AOI21X1 U8440 ( .A0(n9727), .A1(n8348), .B0(n9728), .Y(n9726) );
  AOI21X1 U8441 ( .A0(n8252), .A1(n9729), .B0(n12183), .Y(n9728) );
  NAND3X1 U8442 ( .A(n7926), .B(n9730), .C(n9731), .Y(n9729) );
  INVX1 U8443 ( .A(n9731), .Y(n8348) );
  AOI21X1 U8444 ( .A0(n12299), .A1(n9732), .B0(n9733), .Y(n9731) );
  MX2X1 U8445 ( .A(n9734), .B(n9735), .S0(n7424), .Y(n9733) );
  NAND4X1 U8446 ( .A(n9736), .B(n9737), .C(n9738), .D(n9739), .Y(n9735) );
  OR2X1 U8447 ( .A(n9740), .B(n8255), .Y(n9739) );
  AOI22X1 U8448 ( .A0(n12286), .A1(g17764), .B0(n12285), .B1(g17722), .Y(n9740) );
  AOI22X1 U8449 ( .A0(n9741), .A1(n12297), .B0(n9742), .B1(n12296), .Y(n9738)
         );
  NOR2X1 U8450 ( .A(n5253), .B(n8256), .Y(n9742) );
  INVX1 U8451 ( .A(n9743), .Y(n8256) );
  NOR2X1 U8452 ( .A(n5270), .B(n8258), .Y(n9741) );
  OR2X1 U8453 ( .A(n9744), .B(n8257), .Y(n9737) );
  AOI22X1 U8454 ( .A0(n12293), .A1(g13099), .B0(n12295), .B1(n12294), .Y(n9744) );
  MX2X1 U8455 ( .A(n9745), .B(n9746), .S0(g12470), .Y(n9736) );
  AOI21X1 U8456 ( .A0(n9743), .A1(n7388), .B0(n9747), .Y(n9746) );
  INVX1 U8457 ( .A(n9748), .Y(n9745) );
  NAND4X1 U8458 ( .A(n9749), .B(n9750), .C(n9751), .D(n9752), .Y(n9734) );
  NAND3X1 U8459 ( .A(n9743), .B(g17764), .C(n12284), .Y(n9752) );
  AOI22X1 U8460 ( .A0(n9753), .A1(n12282), .B0(n9754), .B1(n12283), .Y(n9751)
         );
  NOR2X1 U8461 ( .A(n5270), .B(n8257), .Y(n9754) );
  INVX1 U8462 ( .A(n9718), .Y(n8257) );
  NOR2X1 U8463 ( .A(n5253), .B(n8255), .Y(n9753) );
  INVX1 U8464 ( .A(n9755), .Y(n8255) );
  OR2X1 U8465 ( .A(n9756), .B(n8258), .Y(n9750) );
  INVX1 U8466 ( .A(n9757), .Y(n8258) );
  AOI22X1 U8467 ( .A0(n12279), .A1(g13099), .B0(n12280), .B1(n12294), .Y(n9756) );
  MX2X1 U8468 ( .A(n9758), .B(n9759), .S0(g12470), .Y(n9749) );
  AOI21X1 U8469 ( .A0(n9755), .A1(n7441), .B0(n9748), .Y(n9759) );
  NAND3X1 U8470 ( .A(n9760), .B(n9761), .C(n9762), .Y(n9748) );
  NAND3X1 U8471 ( .A(n9743), .B(g17778), .C(n12292), .Y(n9762) );
  NAND3X1 U8472 ( .A(n9718), .B(g14828), .C(n12291), .Y(n9761) );
  NAND3X1 U8473 ( .A(n9757), .B(g17688), .C(n12290), .Y(n9760) );
  INVX1 U8474 ( .A(n9747), .Y(n9758) );
  NAND3X1 U8475 ( .A(n9763), .B(n9764), .C(n9765), .Y(n9747) );
  NAND3X1 U8476 ( .A(n9757), .B(g14828), .C(n12289), .Y(n9765) );
  NOR2X1 U8477 ( .A(n7248), .B(n12305), .Y(n9757) );
  NAND3X1 U8478 ( .A(n9755), .B(g17778), .C(n12287), .Y(n9764) );
  NOR2X1 U8479 ( .A(n12304), .B(n12305), .Y(n9755) );
  NAND3X1 U8480 ( .A(n9718), .B(g17688), .C(n12288), .Y(n9763) );
  NOR2X1 U8481 ( .A(n7248), .B(n7544), .Y(n9718) );
  INVX1 U8482 ( .A(n9730), .Y(n9732) );
  INVX1 U8483 ( .A(n9766), .Y(n9727) );
  AOI21X1 U8484 ( .A0(n8249), .A1(n12183), .B0(n9767), .Y(n9766) );
  AOI22X1 U8485 ( .A0(n12184), .A1(n7898), .B0(n12187), .B1(test_se), .Y(n9725) );
  OAI21X1 U8486 ( .A0(n12183), .A1(n7870), .B0(n9768), .Y(n6554) );
  AOI22X1 U8487 ( .A0(n12180), .A1(n9769), .B0(n9770), .B1(n12184), .Y(n9768)
         );
  OAI21X1 U8488 ( .A0(test_se), .A1(n8556), .B0(n7919), .Y(n9769) );
  INVX1 U8489 ( .A(n9771), .Y(n8556) );
  OAI21X1 U8490 ( .A0(n9772), .A1(n7318), .B0(n9773), .Y(n6553) );
  NOR2X1 U8491 ( .A(n9774), .B(n9775), .Y(n9773) );
  AOI21X1 U8492 ( .A0(n7921), .A1(n9776), .B0(n12183), .Y(n9775) );
  NAND3X1 U8493 ( .A(n7678), .B(n7870), .C(n9777), .Y(n9776) );
  AOI21X1 U8494 ( .A0(n7870), .A1(n9778), .B0(n7678), .Y(n9774) );
  NAND3X1 U8495 ( .A(n12183), .B(g35), .C(n9777), .Y(n9778) );
  OAI21X1 U8496 ( .A0(n9779), .A1(n7567), .B0(n9780), .Y(n6552) );
  MX2X1 U8497 ( .A(n9781), .B(n7318), .S0(n7956), .Y(n9780) );
  NAND2X1 U8498 ( .A(n9771), .B(n7567), .Y(n9781) );
  OAI21X1 U8499 ( .A0(n9772), .A1(n7656), .B0(n9782), .Y(n6551) );
  OAI21X1 U8500 ( .A0(n9777), .A1(n8593), .B0(n12176), .Y(n9782) );
  OAI21X1 U8501 ( .A0(n9772), .A1(n7579), .B0(n9783), .Y(n6550) );
  MX2X1 U8502 ( .A(n9784), .B(n9785), .S0(n7656), .Y(n9783) );
  NAND2X1 U8503 ( .A(n9767), .B(n7567), .Y(n9785) );
  INVX1 U8504 ( .A(n9786), .Y(n9767) );
  AOI21X1 U8505 ( .A0(n12176), .A1(n9777), .B0(n8593), .Y(n9784) );
  OAI21X1 U8506 ( .A0(n7926), .A1(n7579), .B0(n9787), .Y(n6549) );
  MX2X1 U8507 ( .A(n9772), .B(n9786), .S0(n7582), .Y(n9787) );
  NAND2X1 U8508 ( .A(n9777), .B(n7926), .Y(n9786) );
  NOR2X1 U8509 ( .A(n9730), .B(n9721), .Y(n9777) );
  AOI21X1 U8510 ( .A0(n9730), .A1(n7926), .B0(n8349), .Y(n9772) );
  NAND3X1 U8511 ( .A(n9743), .B(g17722), .C(n12298), .Y(n9730) );
  NOR2X1 U8512 ( .A(n7544), .B(n12304), .Y(n9743) );
  MX2X1 U8513 ( .A(n12174), .B(n12175), .S0(n9779), .Y(n6548) );
  OAI21X1 U8514 ( .A0(n7323), .A1(n9779), .B0(n9788), .Y(n6547) );
  MX2X1 U8515 ( .A(n9789), .B(n9790), .S0(n12174), .Y(n9788) );
  AOI21X1 U8516 ( .A0(n12175), .A1(n9771), .B0(n8593), .Y(n9790) );
  NAND3X1 U8517 ( .A(n7926), .B(n7582), .C(n9771), .Y(n9789) );
  INVX1 U8518 ( .A(n9770), .Y(n9779) );
  INVX1 U8519 ( .A(n9791), .Y(n6546) );
  AOI22X1 U8520 ( .A0(n12173), .A1(n9792), .B0(n12180), .B1(test_se), .Y(n9791) );
  NAND2X1 U8521 ( .A(n9793), .B(n9794), .Y(n6545) );
  MX2X1 U8522 ( .A(n9795), .B(n12173), .S0(n7956), .Y(n9793) );
  INVX1 U8523 ( .A(n9796), .Y(n6544) );
  AOI22X1 U8524 ( .A0(n9797), .A1(n7260), .B0(n7955), .B1(n7426), .Y(n9796) );
  OAI21X1 U8525 ( .A0(n12182), .A1(n9798), .B0(n9799), .Y(n6543) );
  OAI21X1 U8526 ( .A0(n12182), .A1(n7962), .B0(n12181), .Y(n9799) );
  INVX1 U8527 ( .A(n9792), .Y(n9798) );
  NAND2X1 U8528 ( .A(n9800), .B(n9801), .Y(n6542) );
  MX2X1 U8529 ( .A(n9802), .B(n12182), .S0(n7957), .Y(n9801) );
  AOI21X1 U8530 ( .A0(n9792), .A1(n12185), .B0(n9803), .Y(n9800) );
  NOR2X1 U8531 ( .A(n7956), .B(n12181), .Y(n9792) );
  OAI21X1 U8532 ( .A0(n8534), .A1(n9804), .B0(n9805), .Y(n6541) );
  MX2X1 U8533 ( .A(n9806), .B(n7482), .S0(n7957), .Y(n9805) );
  NAND2X1 U8534 ( .A(n12279), .B(n9804), .Y(n9806) );
  OR2X1 U8535 ( .A(n9807), .B(n9808), .Y(n9804) );
  NAND2X1 U8536 ( .A(n9809), .B(n9810), .Y(n6540) );
  MX2X1 U8537 ( .A(n9811), .B(n8534), .S0(n9812), .Y(n9810) );
  NOR2X1 U8538 ( .A(n7260), .B(n9802), .Y(n9812) );
  NAND2X1 U8539 ( .A(n12295), .B(n7926), .Y(n9811) );
  AOI22X1 U8540 ( .A0(n12286), .A1(n7896), .B0(test_se), .B1(n7388), .Y(n9809)
         );
  NAND2X1 U8541 ( .A(n9813), .B(n9814), .Y(n6539) );
  MX2X1 U8542 ( .A(n9815), .B(n8534), .S0(n9816), .Y(n9814) );
  NOR2X1 U8543 ( .A(n9807), .B(n9794), .Y(n9816) );
  NAND2X1 U8544 ( .A(n12282), .B(n7926), .Y(n9815) );
  AOI22X1 U8545 ( .A0(n12279), .A1(n7896), .B0(n12295), .B1(test_se), .Y(n9813) );
  NAND2X1 U8546 ( .A(n9817), .B(n9818), .Y(n6538) );
  MX2X1 U8547 ( .A(n9819), .B(n8534), .S0(n9820), .Y(n9818) );
  NOR2X1 U8548 ( .A(n9795), .B(n9807), .Y(n9820) );
  NAND2X1 U8549 ( .A(n12283), .B(n7926), .Y(n9819) );
  AOI22X1 U8550 ( .A0(n12282), .A1(n7896), .B0(n12289), .B1(test_se), .Y(n9817) );
  NAND2X1 U8551 ( .A(n9821), .B(n9822), .Y(n6537) );
  MX2X1 U8552 ( .A(n9823), .B(n8534), .S0(n9824), .Y(n9822) );
  NOR2X1 U8553 ( .A(n9825), .B(n9807), .Y(n9824) );
  NAND2X1 U8554 ( .A(n12284), .B(n7926), .Y(n9823) );
  AOI22X1 U8555 ( .A0(n12283), .A1(n7896), .B0(n12287), .B1(test_se), .Y(n9821) );
  NAND2X1 U8556 ( .A(n9826), .B(n9827), .Y(n6536) );
  MX2X1 U8557 ( .A(n9828), .B(n8534), .S0(n9829), .Y(n9827) );
  NOR2X1 U8558 ( .A(n7260), .B(n9807), .Y(n9829) );
  NAND2X1 U8559 ( .A(n12182), .B(n7482), .Y(n9807) );
  NAND2X1 U8560 ( .A(n12280), .B(n7926), .Y(n9828) );
  AOI22X1 U8561 ( .A0(n12284), .A1(n7896), .B0(test_se), .B1(n7441), .Y(n9826)
         );
  NAND2X1 U8562 ( .A(n9830), .B(n9831), .Y(n6535) );
  AOI22X1 U8563 ( .A0(n9832), .A1(n7926), .B0(n9833), .B1(n9834), .Y(n9831) );
  AOI21X1 U8564 ( .A0(n9834), .A1(n9835), .B0(n12281), .Y(n9832) );
  INVX1 U8565 ( .A(n9808), .Y(n9834) );
  AOI22X1 U8566 ( .A0(n12280), .A1(n7896), .B0(n12279), .B1(test_se), .Y(n9830) );
  NAND2X1 U8567 ( .A(n9836), .B(n9837), .Y(n6534) );
  AOI22X1 U8568 ( .A0(n9838), .A1(n12291), .B0(n9833), .B1(n9839), .Y(n9837)
         );
  AOI21X1 U8569 ( .A0(n9839), .A1(n9835), .B0(n7961), .Y(n9838) );
  AOI22X1 U8570 ( .A0(n7896), .A1(n7441), .B0(n12282), .B1(test_se), .Y(n9836)
         );
  NAND2X1 U8571 ( .A(n9840), .B(n9841), .Y(n6533) );
  AOI22X1 U8572 ( .A0(n9842), .A1(n12292), .B0(n9833), .B1(n9843), .Y(n9841)
         );
  AOI21X1 U8573 ( .A0(n9835), .A1(n9843), .B0(n7958), .Y(n9842) );
  INVX1 U8574 ( .A(n9795), .Y(n9843) );
  AOI22X1 U8575 ( .A0(n12291), .A1(n7896), .B0(n12283), .B1(test_se), .Y(n9840) );
  NAND2X1 U8576 ( .A(n9844), .B(n9845), .Y(n6532) );
  AOI22X1 U8577 ( .A0(n9846), .A1(n12290), .B0(n9833), .B1(n9797), .Y(n9845)
         );
  AOI21X1 U8578 ( .A0(n9835), .A1(n9797), .B0(n7963), .Y(n9846) );
  AOI22X1 U8579 ( .A0(n12292), .A1(n7896), .B0(n12284), .B1(test_se), .Y(n9844) );
  NAND2X1 U8580 ( .A(n9847), .B(n9848), .Y(n6531) );
  AOI22X1 U8581 ( .A0(n9849), .A1(n12285), .B0(n9833), .B1(n12181), .Y(n9848)
         );
  AND2X1 U8582 ( .A(n9835), .B(n8893), .Y(n9833) );
  NOR2X1 U8583 ( .A(n9803), .B(n7961), .Y(n9849) );
  AND2X1 U8584 ( .A(n9835), .B(n12181), .Y(n9803) );
  NOR2X1 U8585 ( .A(n12185), .B(n12182), .Y(n9835) );
  AOI22X1 U8586 ( .A0(n12290), .A1(n7896), .B0(n12293), .B1(test_se), .Y(n9847) );
  NAND2X1 U8587 ( .A(n9850), .B(n9851), .Y(n6530) );
  MX2X1 U8588 ( .A(n9852), .B(n8534), .S0(n9853), .Y(n9851) );
  NOR2X1 U8589 ( .A(n9802), .B(n9808), .Y(n9853) );
  NAND2X1 U8590 ( .A(n12293), .B(n7927), .Y(n9852) );
  AOI22X1 U8591 ( .A0(n12285), .A1(n7896), .B0(n12280), .B1(test_se), .Y(n9850) );
  NAND2X1 U8592 ( .A(n9854), .B(n9855), .Y(n6529) );
  MX2X1 U8593 ( .A(n9856), .B(n8534), .S0(n9857), .Y(n9855) );
  NOR2X1 U8594 ( .A(n9802), .B(n9794), .Y(n9857) );
  NAND2X1 U8595 ( .A(n12296), .B(n7927), .Y(n9856) );
  AOI22X1 U8596 ( .A0(n12293), .A1(n7896), .B0(n12291), .B1(test_se), .Y(n9854) );
  NAND2X1 U8597 ( .A(n9858), .B(n9859), .Y(n6528) );
  MX2X1 U8598 ( .A(n9860), .B(n8534), .S0(n9861), .Y(n9859) );
  NOR2X1 U8599 ( .A(n9795), .B(n9802), .Y(n9861) );
  NAND2X1 U8600 ( .A(n12297), .B(n7927), .Y(n9860) );
  AOI22X1 U8601 ( .A0(n12296), .A1(n7895), .B0(n12292), .B1(test_se), .Y(n9858) );
  NAND2X1 U8602 ( .A(n9862), .B(n9863), .Y(n6527) );
  MX2X1 U8603 ( .A(n9864), .B(n8534), .S0(n9865), .Y(n9863) );
  NOR2X1 U8604 ( .A(n9866), .B(n9808), .Y(n9865) );
  NAND3X1 U8605 ( .A(n12173), .B(n7260), .C(n12172), .Y(n9808) );
  NAND2X1 U8606 ( .A(n7927), .B(n7388), .Y(n9864) );
  AOI22X1 U8607 ( .A0(n12295), .A1(n7895), .B0(n12285), .B1(test_se), .Y(n9862) );
  NAND2X1 U8608 ( .A(n9867), .B(n9868), .Y(n6526) );
  MX2X1 U8609 ( .A(n9869), .B(n8534), .S0(n9870), .Y(n9868) );
  NOR2X1 U8610 ( .A(n9866), .B(n9794), .Y(n9870) );
  INVX1 U8611 ( .A(n9839), .Y(n9794) );
  NOR2X1 U8612 ( .A(n7426), .B(n12173), .Y(n9839) );
  NAND2X1 U8613 ( .A(n12289), .B(n7927), .Y(n9869) );
  AOI22X1 U8614 ( .A0(n7895), .A1(n7388), .B0(n12296), .B1(test_se), .Y(n9867)
         );
  NAND2X1 U8615 ( .A(n9871), .B(n9872), .Y(n6525) );
  MX2X1 U8616 ( .A(n9873), .B(n8534), .S0(n9874), .Y(n9872) );
  NOR2X1 U8617 ( .A(n9866), .B(n9795), .Y(n9874) );
  NAND2X1 U8618 ( .A(n12173), .B(n7426), .Y(n9795) );
  NAND2X1 U8619 ( .A(n12287), .B(n7927), .Y(n9873) );
  AOI22X1 U8620 ( .A0(n12289), .A1(n7895), .B0(n12297), .B1(test_se), .Y(n9871) );
  NAND2X1 U8621 ( .A(n9875), .B(n9876), .Y(n6524) );
  MX2X1 U8622 ( .A(n9877), .B(n8534), .S0(n9878), .Y(n9876) );
  NOR2X1 U8623 ( .A(n9825), .B(n9802), .Y(n9878) );
  NAND2X1 U8624 ( .A(n12182), .B(n12185), .Y(n9802) );
  NAND2X1 U8625 ( .A(n12286), .B(n7927), .Y(n9877) );
  AOI22X1 U8626 ( .A0(n12297), .A1(n7895), .B0(n12290), .B1(test_se), .Y(n9875) );
  NAND2X1 U8627 ( .A(n9879), .B(n9880), .Y(n6523) );
  MX2X1 U8628 ( .A(n9881), .B(n8534), .S0(n9882), .Y(n9880) );
  NOR2X1 U8629 ( .A(n9866), .B(n9825), .Y(n9882) );
  INVX1 U8630 ( .A(n9797), .Y(n9825) );
  NOR2X1 U8631 ( .A(n12173), .B(n12172), .Y(n9797) );
  NAND2X1 U8632 ( .A(n12288), .B(n7927), .Y(n9881) );
  AOI22X1 U8633 ( .A0(n12287), .A1(n7895), .B0(n12286), .B1(test_se), .Y(n9879) );
  OAI21X1 U8634 ( .A0(n7927), .A1(n7796), .B0(n9883), .Y(n6522) );
  AOI22X1 U8635 ( .A0(n9770), .A1(n12299), .B0(n9771), .B1(n8893), .Y(n9883)
         );
  NOR2X1 U8636 ( .A(n7961), .B(n9771), .Y(n9770) );
  NOR2X1 U8637 ( .A(n7260), .B(n9866), .Y(n9771) );
  OR2X1 U8638 ( .A(n7482), .B(n12182), .Y(n9866) );
  NAND2X1 U8639 ( .A(n9884), .B(n9885), .Y(n6521) );
  MX2X1 U8640 ( .A(n9886), .B(n9887), .S0(n7376), .Y(n9885) );
  NAND2X1 U8641 ( .A(n9888), .B(n7927), .Y(n9887) );
  OR2X1 U8642 ( .A(n9889), .B(n9888), .Y(n9886) );
  NOR2X1 U8643 ( .A(n12277), .B(n12278), .Y(n9888) );
  AOI22X1 U8644 ( .A0(n12278), .A1(n7895), .B0(n12387), .B1(test_se), .Y(n9884) );
  NAND2X1 U8645 ( .A(n9890), .B(n9891), .Y(n6520) );
  MX2X1 U8646 ( .A(n9892), .B(n7870), .S0(n12278), .Y(n9891) );
  NAND3X1 U8647 ( .A(n9893), .B(n7270), .C(n12276), .Y(n9892) );
  AOI22X1 U8648 ( .A0(n9894), .A1(n7927), .B0(n9895), .B1(n7376), .Y(n9890) );
  OAI21X1 U8649 ( .A0(test_se), .A1(n9896), .B0(n7919), .Y(n9895) );
  MX2X1 U8650 ( .A(n7270), .B(n9897), .S0(n7406), .Y(n9896) );
  NAND2X1 U8651 ( .A(n9898), .B(n7270), .Y(n9897) );
  OAI21X1 U8652 ( .A0(n12271), .A1(n7927), .B0(n9899), .Y(n6519) );
  MX2X1 U8653 ( .A(n9900), .B(n9901), .S0(n7399), .Y(n9899) );
  AOI21X1 U8654 ( .A0(n9894), .A1(n7927), .B0(n9902), .Y(n9901) );
  NAND3X1 U8655 ( .A(n9903), .B(n9904), .C(n9893), .Y(n9900) );
  OAI21X1 U8656 ( .A0(n7962), .A1(n9905), .B0(n9906), .Y(n6518) );
  AOI22X1 U8657 ( .A0(n9907), .A1(n9908), .B0(n12270), .B1(n9909), .Y(n9906)
         );
  OAI21X1 U8658 ( .A0(n9903), .A1(n7427), .B0(n7922), .Y(n9909) );
  MX2X1 U8659 ( .A(n9903), .B(n9904), .S0(n7399), .Y(n9908) );
  NOR2X1 U8660 ( .A(n12269), .B(n9889), .Y(n9907) );
  NAND2X1 U8661 ( .A(n9910), .B(n9911), .Y(n6517) );
  MX2X1 U8662 ( .A(n12268), .B(n9912), .S0(n9913), .Y(n9911) );
  NAND3X1 U8663 ( .A(n9893), .B(n9905), .C(n12268), .Y(n9912) );
  AOI21X1 U8664 ( .A0(n7961), .A1(n7427), .B0(n9914), .Y(n9910) );
  INVX1 U8665 ( .A(n9915), .Y(n9914) );
  NAND2X1 U8666 ( .A(n9916), .B(n9917), .Y(n6516) );
  MX2X1 U8667 ( .A(n9918), .B(n9919), .S0(n7408), .Y(n9916) );
  NAND3X1 U8668 ( .A(n9905), .B(n7358), .C(n9893), .Y(n9919) );
  NOR2X1 U8669 ( .A(n7962), .B(n9920), .Y(n9918) );
  MX2X1 U8670 ( .A(n9921), .B(n9922), .S0(n7358), .Y(n9920) );
  NOR2X1 U8671 ( .A(n9921), .B(n9889), .Y(n9922) );
  NAND2X1 U8672 ( .A(n9923), .B(n9924), .Y(n6515) );
  MX2X1 U8673 ( .A(n9925), .B(n8721), .S0(n7358), .Y(n9924) );
  NAND2X1 U8674 ( .A(n9926), .B(n9893), .Y(n9925) );
  AOI21X1 U8675 ( .A0(n9927), .A1(n7408), .B0(n12273), .Y(n9926) );
  AOI22X1 U8676 ( .A0(n9928), .A1(n9898), .B0(n12273), .B1(n9929), .Y(n9923)
         );
  OAI21X1 U8677 ( .A0(n12274), .A1(n9930), .B0(n9917), .Y(n9929) );
  INVX1 U8678 ( .A(n9931), .Y(n9917) );
  AND2X1 U8679 ( .A(n9930), .B(n9932), .Y(n9928) );
  NAND2X1 U8680 ( .A(n12268), .B(n9921), .Y(n9930) );
  OAI21X1 U8681 ( .A0(n12273), .A1(n7927), .B0(n9933), .Y(n6514) );
  MX2X1 U8682 ( .A(n9934), .B(n9935), .S0(n12275), .Y(n9933) );
  AOI21X1 U8683 ( .A0(n9931), .A1(n12273), .B0(n9936), .Y(n9935) );
  INVX1 U8684 ( .A(n9937), .Y(n9936) );
  NOR2X1 U8685 ( .A(n9915), .B(n7358), .Y(n9931) );
  NAND3X1 U8686 ( .A(n7927), .B(n7408), .C(n9927), .Y(n9915) );
  INVX1 U8687 ( .A(n9905), .Y(n9927) );
  NAND3X1 U8688 ( .A(n9894), .B(n7399), .C(n12269), .Y(n9905) );
  INVX1 U8689 ( .A(n9904), .Y(n9894) );
  NAND3X1 U8690 ( .A(n12276), .B(n12278), .C(n12271), .Y(n9904) );
  NAND2X1 U8691 ( .A(n9893), .B(n9937), .Y(n9934) );
  NAND3X1 U8692 ( .A(n9921), .B(n9932), .C(n12268), .Y(n9937) );
  INVX1 U8693 ( .A(n9913), .Y(n9921) );
  NAND3X1 U8694 ( .A(n12270), .B(n7427), .C(n9902), .Y(n9913) );
  INVX1 U8695 ( .A(n9903), .Y(n9902) );
  NAND3X1 U8696 ( .A(n7376), .B(n7270), .C(n12277), .Y(n9903) );
  INVX1 U8697 ( .A(n9889), .Y(n9893) );
  NAND2X1 U8698 ( .A(n9898), .B(n7927), .Y(n9889) );
  MX2X1 U8699 ( .A(n9938), .B(n9939), .S0(n12275), .Y(n9898) );
  NAND2X1 U8700 ( .A(n12277), .B(n9932), .Y(n9939) );
  OAI21X1 U8701 ( .A0(n12275), .A1(n7870), .B0(n9940), .Y(n6513) );
  AOI22X1 U8702 ( .A0(n9941), .A1(n3816), .B0(n12266), .B1(n7895), .Y(n9940)
         );
  NOR2X1 U8703 ( .A(n9942), .B(n7962), .Y(n9941) );
  AOI21X1 U8704 ( .A0(g9497), .A1(n7797), .B0(n12277), .Y(n9942) );
  OAI21X1 U8705 ( .A0(n7869), .A1(n7406), .B0(n9943), .Y(n6512) );
  MX2X1 U8706 ( .A(n9944), .B(n7962), .S0(n12275), .Y(n9943) );
  AOI21X1 U8707 ( .A0(n9938), .A1(n7869), .B0(n7895), .Y(n9944) );
  NAND3X1 U8708 ( .A(n12274), .B(n12278), .C(n12273), .Y(n9938) );
  MX2X1 U8709 ( .A(n9945), .B(n12265), .S0(n7958), .Y(n6511) );
  NAND3X1 U8710 ( .A(n12277), .B(n9932), .C(n12275), .Y(n9945) );
  NOR2X1 U8711 ( .A(n12274), .B(n12273), .Y(n9932) );
  AOI21X1 U8712 ( .A0(n8721), .A1(n7349), .B0(n7750), .Y(n6510) );
  NAND2X1 U8713 ( .A(n9946), .B(n9947), .Y(n6509) );
  NAND3X1 U8714 ( .A(n7750), .B(n7327), .C(n7927), .Y(n9947) );
  MX2X1 U8715 ( .A(n9948), .B(n9949), .S0(n12262), .Y(n9946) );
  OAI21X1 U8716 ( .A0(n12265), .A1(n12263), .B0(n9948), .Y(n9949) );
  AOI21X1 U8717 ( .A0(n9950), .A1(n7927), .B0(n12263), .Y(n6508) );
  MX2X1 U8718 ( .A(n12264), .B(n12265), .S0(n7243), .Y(n9950) );
  OAI21X1 U8719 ( .A0(n9951), .A1(n7471), .B0(n9952), .Y(n6507) );
  OAI21X1 U8720 ( .A0(n8593), .A1(n7471), .B0(n7243), .Y(n9952) );
  INVX1 U8721 ( .A(n9948), .Y(n9951) );
  OAI22X1 U8722 ( .A0(n12260), .A1(n9953), .B0(n9954), .B1(n7471), .Y(n6506)
         );
  AOI21X1 U8723 ( .A0(n12260), .A1(n7243), .B0(n7962), .Y(n9954) );
  AOI21X1 U8724 ( .A0(n7927), .A1(n7471), .B0(n9948), .Y(n9953) );
  INVX1 U8725 ( .A(n9955), .Y(n6505) );
  AOI22X1 U8726 ( .A0(n12259), .A1(n7927), .B0(test_se), .B1(n7498), .Y(n9955)
         );
  OAI21X1 U8727 ( .A0(n3814), .A1(n7869), .B0(n9956), .Y(n6504) );
  AOI21X1 U8728 ( .A0(n12277), .A1(n7895), .B0(n9957), .Y(n9956) );
  NAND2X1 U8729 ( .A(n9958), .B(n9959), .Y(n6503) );
  AOI21X1 U8730 ( .A0(n9960), .A1(n9961), .B0(n9962), .Y(n9959) );
  AOI21X1 U8731 ( .A0(n9963), .A1(n9964), .B0(n12257), .Y(n9962) );
  NAND3X1 U8732 ( .A(n9965), .B(n9966), .C(n7927), .Y(n9964) );
  INVX1 U8733 ( .A(n9960), .Y(n9965) );
  INVX1 U8734 ( .A(n9967), .Y(n9961) );
  AOI21X1 U8735 ( .A0(n9968), .A1(n12257), .B0(n9969), .Y(n9967) );
  AOI22X1 U8736 ( .A0(n12258), .A1(n7895), .B0(n12272), .B1(test_se), .Y(n9958) );
  OAI21X1 U8737 ( .A0(n12257), .A1(n7921), .B0(n9970), .Y(n6502) );
  AOI21X1 U8738 ( .A0(n9971), .A1(n7869), .B0(n9972), .Y(n9970) );
  AOI21X1 U8739 ( .A0(n7869), .A1(n9973), .B0(n7713), .Y(n9972) );
  NAND3X1 U8740 ( .A(n12257), .B(g35), .C(n9974), .Y(n9973) );
  MX2X1 U8741 ( .A(n9975), .B(n9976), .S0(n9974), .Y(n9971) );
  NOR2X1 U8742 ( .A(n12257), .B(n12258), .Y(n9976) );
  OAI21X1 U8743 ( .A0(n9977), .A1(n7568), .B0(n9978), .Y(n6501) );
  MX2X1 U8744 ( .A(n9979), .B(n7823), .S0(n7957), .Y(n9978) );
  NAND2X1 U8745 ( .A(g32975), .B(n7568), .Y(n9979) );
  OAI21X1 U8746 ( .A0(n12252), .A1(n9980), .B0(n9981), .Y(n6500) );
  OAI21X1 U8747 ( .A0(n9974), .A1(n8593), .B0(n12253), .Y(n9981) );
  OAI21X1 U8748 ( .A0(n12694), .A1(n9980), .B0(n9982), .Y(n6499) );
  MX2X1 U8749 ( .A(n9983), .B(n9984), .S0(n12252), .Y(n9982) );
  NAND2X1 U8750 ( .A(n9969), .B(n7568), .Y(n9984) );
  INVX1 U8751 ( .A(n9985), .Y(n9969) );
  AOI21X1 U8752 ( .A0(n12253), .A1(n9974), .B0(n8593), .Y(n9983) );
  OAI21X1 U8753 ( .A0(n12694), .A1(n7927), .B0(n9986), .Y(n6498) );
  MX2X1 U8754 ( .A(n9980), .B(n9985), .S0(n7583), .Y(n9986) );
  NAND2X1 U8755 ( .A(n9974), .B(n7927), .Y(n9985) );
  OR2X1 U8756 ( .A(n7963), .B(n9974), .Y(n9980) );
  NOR2X1 U8757 ( .A(n9966), .B(n9987), .Y(n9974) );
  NAND3X1 U8758 ( .A(g25219), .B(g17577), .C(g25114), .Y(n9966) );
  MX2X1 U8759 ( .A(n12250), .B(n12251), .S0(n9977), .Y(n6497) );
  OAI21X1 U8760 ( .A0(n9977), .A1(n7646), .B0(n9988), .Y(n6496) );
  MX2X1 U8761 ( .A(n9989), .B(n9990), .S0(n12250), .Y(n9988) );
  AOI21X1 U8762 ( .A0(n12251), .A1(g32975), .B0(n8593), .Y(n9990) );
  NAND3X1 U8763 ( .A(n7927), .B(n7583), .C(g32975), .Y(n9989) );
  INVX1 U8764 ( .A(n8496), .Y(n9977) );
  INVX1 U8765 ( .A(n9991), .Y(n6495) );
  AOI22X1 U8766 ( .A0(n12249), .A1(n9992), .B0(n12254), .B1(test_se), .Y(n9991) );
  NAND2X1 U8767 ( .A(n9993), .B(n9994), .Y(n6494) );
  MX2X1 U8768 ( .A(n9995), .B(n12249), .S0(n7956), .Y(n9993) );
  INVX1 U8769 ( .A(n9996), .Y(n6493) );
  AOI22X1 U8770 ( .A0(n9997), .A1(n7264), .B0(n7963), .B1(n7428), .Y(n9996) );
  OAI21X1 U8771 ( .A0(n12256), .A1(n9998), .B0(n9999), .Y(n6492) );
  OAI21X1 U8772 ( .A0(n12256), .A1(n7963), .B0(n12255), .Y(n9999) );
  INVX1 U8773 ( .A(n9992), .Y(n9998) );
  NAND2X1 U8774 ( .A(n10000), .B(n10001), .Y(n6491) );
  MX2X1 U8775 ( .A(n10002), .B(n12256), .S0(n7961), .Y(n10001) );
  AOI21X1 U8776 ( .A0(n9992), .A1(n12259), .B0(n10003), .Y(n10000) );
  NOR2X1 U8777 ( .A(n7963), .B(n12255), .Y(n9992) );
  OAI21X1 U8778 ( .A0(n8534), .A1(n10004), .B0(n10005), .Y(n6490) );
  MX2X1 U8779 ( .A(n10006), .B(n7493), .S0(n7955), .Y(n10005) );
  NAND2X1 U8780 ( .A(n12975), .B(n10004), .Y(n10006) );
  OR2X1 U8781 ( .A(n10007), .B(n10008), .Y(n10004) );
  NAND2X1 U8782 ( .A(n10009), .B(n10010), .Y(n6489) );
  MX2X1 U8783 ( .A(n10011), .B(n8534), .S0(n10012), .Y(n10010) );
  NOR2X1 U8784 ( .A(n7264), .B(n10002), .Y(n10012) );
  NAND2X1 U8785 ( .A(n12981), .B(n7928), .Y(n10011) );
  AOI22X1 U8786 ( .A0(n12990), .A1(n7895), .B0(n12985), .B1(test_se), .Y(
        n10009) );
  NAND2X1 U8787 ( .A(n10013), .B(n10014), .Y(n6488) );
  MX2X1 U8788 ( .A(n10015), .B(n8534), .S0(n10016), .Y(n10014) );
  NOR2X1 U8789 ( .A(n10007), .B(n9994), .Y(n10016) );
  NAND2X1 U8790 ( .A(n12977), .B(n7928), .Y(n10015) );
  AOI22X1 U8791 ( .A0(n12975), .A1(n7894), .B0(n12981), .B1(test_se), .Y(
        n10013) );
  NAND2X1 U8792 ( .A(n10017), .B(n10018), .Y(n6487) );
  MX2X1 U8793 ( .A(n10019), .B(n8534), .S0(n10020), .Y(n10018) );
  NOR2X1 U8794 ( .A(n9995), .B(n10007), .Y(n10020) );
  NAND2X1 U8795 ( .A(n12978), .B(n7928), .Y(n10019) );
  AOI22X1 U8796 ( .A0(n12977), .A1(n7894), .B0(n12982), .B1(test_se), .Y(
        n10017) );
  NAND2X1 U8797 ( .A(n10021), .B(n10022), .Y(n6486) );
  MX2X1 U8798 ( .A(n10023), .B(n8534), .S0(n10024), .Y(n10022) );
  NOR2X1 U8799 ( .A(n10025), .B(n10007), .Y(n10024) );
  NAND2X1 U8800 ( .A(n7928), .B(n7227), .Y(n10023) );
  AOI22X1 U8801 ( .A0(n12978), .A1(n7894), .B0(n12983), .B1(test_se), .Y(
        n10021) );
  NAND2X1 U8802 ( .A(n10026), .B(n10027), .Y(n6485) );
  MX2X1 U8803 ( .A(n10028), .B(n8534), .S0(n10029), .Y(n10027) );
  NOR2X1 U8804 ( .A(n7264), .B(n10007), .Y(n10029) );
  NAND2X1 U8805 ( .A(n12256), .B(n7493), .Y(n10007) );
  NAND2X1 U8806 ( .A(n12976), .B(n7928), .Y(n10028) );
  AOI22X1 U8807 ( .A0(n7894), .A1(n7227), .B0(test_se), .B1(n7446), .Y(n10026)
         );
  NAND2X1 U8808 ( .A(n10030), .B(n10031), .Y(n6484) );
  AOI22X1 U8809 ( .A0(n10032), .A1(n7928), .B0(n10033), .B1(n10034), .Y(n10031) );
  AOI21X1 U8810 ( .A0(n10034), .A1(n10035), .B0(n12974), .Y(n10032) );
  INVX1 U8811 ( .A(n10008), .Y(n10034) );
  AOI22X1 U8812 ( .A0(n12976), .A1(n7894), .B0(n12975), .B1(test_se), .Y(
        n10030) );
  NAND2X1 U8813 ( .A(n10036), .B(n10037), .Y(n6483) );
  AOI22X1 U8814 ( .A0(n10038), .A1(n12987), .B0(n10033), .B1(n10039), .Y(
        n10037) );
  AOI21X1 U8815 ( .A0(n10039), .A1(n10035), .B0(n7963), .Y(n10038) );
  AOI22X1 U8816 ( .A0(n7894), .A1(n7446), .B0(n12977), .B1(test_se), .Y(n10036) );
  NAND2X1 U8817 ( .A(n10040), .B(n10041), .Y(n6482) );
  AOI22X1 U8818 ( .A0(n10042), .A1(n12986), .B0(n10033), .B1(n10043), .Y(
        n10041) );
  AOI21X1 U8819 ( .A0(n10035), .A1(n10043), .B0(n7963), .Y(n10042) );
  INVX1 U8820 ( .A(n9995), .Y(n10043) );
  AOI22X1 U8821 ( .A0(n12987), .A1(n7894), .B0(n12978), .B1(test_se), .Y(
        n10040) );
  NAND2X1 U8822 ( .A(n10044), .B(n10045), .Y(n6481) );
  AOI22X1 U8823 ( .A0(n10046), .A1(n12988), .B0(n10033), .B1(n9997), .Y(n10045) );
  AOI21X1 U8824 ( .A0(n10035), .A1(n9997), .B0(n7950), .Y(n10046) );
  AOI22X1 U8825 ( .A0(n12986), .A1(n7894), .B0(test_se), .B1(n7227), .Y(n10044) );
  NAND2X1 U8826 ( .A(n10047), .B(n10048), .Y(n6480) );
  AOI22X1 U8827 ( .A0(n10049), .A1(n12989), .B0(n10033), .B1(n12255), .Y(
        n10048) );
  AND2X1 U8828 ( .A(n10035), .B(n8893), .Y(n10033) );
  NOR2X1 U8829 ( .A(n10003), .B(n7953), .Y(n10049) );
  AND2X1 U8830 ( .A(n10035), .B(n12255), .Y(n10003) );
  NOR2X1 U8831 ( .A(n12259), .B(n12256), .Y(n10035) );
  AOI22X1 U8832 ( .A0(n12988), .A1(n7894), .B0(n12979), .B1(test_se), .Y(
        n10047) );
  NAND2X1 U8833 ( .A(n10050), .B(n10051), .Y(n6479) );
  MX2X1 U8834 ( .A(n10052), .B(n8534), .S0(n10053), .Y(n10051) );
  NOR2X1 U8835 ( .A(n10002), .B(n10008), .Y(n10053) );
  NAND2X1 U8836 ( .A(n12979), .B(n7928), .Y(n10052) );
  AOI22X1 U8837 ( .A0(n12989), .A1(n7894), .B0(n12976), .B1(test_se), .Y(
        n10050) );
  NAND2X1 U8838 ( .A(n10054), .B(n10055), .Y(n6478) );
  MX2X1 U8839 ( .A(n10056), .B(n8534), .S0(n10057), .Y(n10055) );
  NOR2X1 U8840 ( .A(n10002), .B(n9994), .Y(n10057) );
  NAND2X1 U8841 ( .A(n12994), .B(n7928), .Y(n10056) );
  AOI22X1 U8842 ( .A0(n12979), .A1(n7894), .B0(n12987), .B1(test_se), .Y(
        n10054) );
  NAND2X1 U8843 ( .A(n10058), .B(n10059), .Y(n6477) );
  MX2X1 U8844 ( .A(n10060), .B(n8534), .S0(n10061), .Y(n10059) );
  NOR2X1 U8845 ( .A(n9995), .B(n10002), .Y(n10061) );
  NAND2X1 U8846 ( .A(n12991), .B(n7928), .Y(n10060) );
  AOI22X1 U8847 ( .A0(n12994), .A1(n7894), .B0(n12986), .B1(test_se), .Y(
        n10058) );
  NAND2X1 U8848 ( .A(n10062), .B(n10063), .Y(n6476) );
  MX2X1 U8849 ( .A(n10064), .B(n8534), .S0(n10065), .Y(n10063) );
  NOR2X1 U8850 ( .A(n10066), .B(n10008), .Y(n10065) );
  NAND3X1 U8851 ( .A(n12249), .B(n7264), .C(n12248), .Y(n10008) );
  NAND2X1 U8852 ( .A(n12985), .B(n7928), .Y(n10064) );
  AOI22X1 U8853 ( .A0(n12981), .A1(n7893), .B0(n12989), .B1(test_se), .Y(
        n10062) );
  NAND2X1 U8854 ( .A(n10067), .B(n10068), .Y(n6475) );
  MX2X1 U8855 ( .A(n10069), .B(n8534), .S0(n10070), .Y(n10068) );
  NOR2X1 U8856 ( .A(n10066), .B(n9994), .Y(n10070) );
  INVX1 U8857 ( .A(n10039), .Y(n9994) );
  NOR2X1 U8858 ( .A(n7428), .B(n12249), .Y(n10039) );
  NAND2X1 U8859 ( .A(n12982), .B(n7928), .Y(n10069) );
  AOI22X1 U8860 ( .A0(n12985), .A1(n7893), .B0(n12994), .B1(test_se), .Y(
        n10067) );
  NAND2X1 U8861 ( .A(n10071), .B(n10072), .Y(n6474) );
  MX2X1 U8862 ( .A(n10073), .B(n8534), .S0(n10074), .Y(n10072) );
  NOR2X1 U8863 ( .A(n10066), .B(n9995), .Y(n10074) );
  NAND2X1 U8864 ( .A(n12249), .B(n7428), .Y(n9995) );
  NAND2X1 U8865 ( .A(n12983), .B(n7928), .Y(n10073) );
  AOI22X1 U8866 ( .A0(n12982), .A1(n7893), .B0(n12991), .B1(test_se), .Y(
        n10071) );
  NAND2X1 U8867 ( .A(n10075), .B(n10076), .Y(n6473) );
  MX2X1 U8868 ( .A(n10077), .B(n8534), .S0(n10078), .Y(n10076) );
  NOR2X1 U8869 ( .A(n10025), .B(n10002), .Y(n10078) );
  NAND2X1 U8870 ( .A(n12256), .B(n12259), .Y(n10002) );
  NAND2X1 U8871 ( .A(n12990), .B(n7928), .Y(n10077) );
  AOI22X1 U8872 ( .A0(n12991), .A1(n7893), .B0(n12988), .B1(test_se), .Y(
        n10075) );
  NAND2X1 U8873 ( .A(n10079), .B(n10080), .Y(n6472) );
  MX2X1 U8874 ( .A(n10081), .B(n8534), .S0(n10082), .Y(n10080) );
  NOR2X1 U8875 ( .A(n10066), .B(n10025), .Y(n10082) );
  INVX1 U8876 ( .A(n9997), .Y(n10025) );
  NOR2X1 U8877 ( .A(n12249), .B(n12248), .Y(n9997) );
  NAND2X1 U8878 ( .A(n12984), .B(n7942), .Y(n10081) );
  AOI22X1 U8879 ( .A0(n12983), .A1(n7893), .B0(n12990), .B1(test_se), .Y(
        n10079) );
  OAI21X1 U8880 ( .A0(n7940), .A1(n7798), .B0(n10083), .Y(n6471) );
  AOI22X1 U8881 ( .A0(n13005), .A1(n8496), .B0(n8893), .B1(g32975), .Y(n10083)
         );
  NOR2X1 U8882 ( .A(n7952), .B(g32975), .Y(n8496) );
  MX2X1 U8883 ( .A(n13005), .B(g17674), .S0(n7849), .Y(n6470) );
  INVX1 U8884 ( .A(n10084), .Y(n6469) );
  MX2X1 U8885 ( .A(n10085), .B(n7869), .S0(g13039), .Y(n10084) );
  NAND4X1 U8886 ( .A(n7821), .B(n5604), .C(n10086), .D(n7940), .Y(n10085) );
  MX2X1 U8887 ( .A(n5605), .B(g12238), .S0(g14662), .Y(n10086) );
  MX2X1 U8888 ( .A(g17577), .B(g12238), .S0(n7848), .Y(n6468) );
  MX2X1 U8889 ( .A(g12238), .B(g14662), .S0(n7848), .Y(n6467) );
  OAI21X1 U8890 ( .A0(n10087), .A1(n10088), .B0(n10089), .Y(n6465) );
  MX2X1 U8891 ( .A(n10090), .B(n7799), .S0(n7961), .Y(n10089) );
  NAND2X1 U8892 ( .A(n10087), .B(n302), .Y(n10090) );
  INVX1 U8893 ( .A(n10091), .Y(n10087) );
  NOR2X1 U8894 ( .A(n10092), .B(n10093), .Y(n6464) );
  MX2X1 U8895 ( .A(n12384), .B(n302), .S0(n7960), .Y(n10093) );
  NOR2X1 U8896 ( .A(n10092), .B(n7657), .Y(n6463) );
  NOR2X1 U8897 ( .A(n10088), .B(n10091), .Y(n10092) );
  NAND4X1 U8898 ( .A(g14662), .B(g17519), .C(g17674), .D(g12238), .Y(n10091)
         );
  INVX1 U8899 ( .A(n9957), .Y(n10088) );
  NOR2X1 U8900 ( .A(n7948), .B(n302), .Y(n9957) );
  OAI21X1 U8901 ( .A0(n7940), .A1(n7626), .B0(n10094), .Y(n6462) );
  MX2X1 U8902 ( .A(n10095), .B(n9963), .S0(n7366), .Y(n10094) );
  INVX1 U8903 ( .A(n10096), .Y(n6461) );
  AOI22X1 U8904 ( .A0(n12240), .A1(n7940), .B0(n12244), .B1(test_se), .Y(
        n10096) );
  OAI21X1 U8905 ( .A0(n7990), .A1(n7869), .B0(n10097), .Y(n6460) );
  AOI21X1 U8906 ( .A0(n12244), .A1(n7893), .B0(n9143), .Y(n10097) );
  NOR2X1 U8907 ( .A(n7954), .B(n12356), .Y(n9143) );
  NAND2X1 U8908 ( .A(n10098), .B(n10099), .Y(n6459) );
  AOI22X1 U8909 ( .A0(n10100), .A1(n12993), .B0(n10101), .B1(n7940), .Y(n10099) );
  AOI21X1 U8910 ( .A0(n7893), .A1(n7366), .B0(n10102), .Y(n10098) );
  MX2X1 U8911 ( .A(g14662), .B(n10103), .S0(n7848), .Y(n10102) );
  NOR2X1 U8912 ( .A(n9987), .B(n10104), .Y(n10103) );
  OAI21X1 U8913 ( .A0(n7869), .A1(n7714), .B0(n10105), .Y(n6458) );
  AOI22X1 U8914 ( .A0(n10106), .A1(n10107), .B0(n10108), .B1(n7459), .Y(n10105) );
  OAI21X1 U8915 ( .A0(n7947), .A1(n10109), .B0(n9963), .Y(n10108) );
  INVX1 U8916 ( .A(n10100), .Y(n9963) );
  AOI21X1 U8917 ( .A0(n10110), .A1(n10111), .B0(n10095), .Y(n10106) );
  INVX1 U8918 ( .A(n9968), .Y(n10095) );
  MX2X1 U8919 ( .A(n10112), .B(n10113), .S0(n7657), .Y(n10111) );
  MX2X1 U8920 ( .A(n10114), .B(n10104), .S0(n7626), .Y(n10110) );
  NAND2X1 U8921 ( .A(n10115), .B(n10116), .Y(n6457) );
  AOI22X1 U8922 ( .A0(n10117), .A1(n7380), .B0(n8345), .B1(n7940), .Y(n10116)
         );
  AOI21X1 U8923 ( .A0(n7893), .A1(n7249), .B0(n10118), .Y(n10115) );
  MX2X1 U8924 ( .A(n7459), .B(n10119), .S0(n7848), .Y(n10118) );
  NOR2X1 U8925 ( .A(n8585), .B(n10120), .Y(n10119) );
  INVX1 U8926 ( .A(n8631), .Y(n8585) );
  INVX1 U8927 ( .A(n10121), .Y(n6456) );
  AOI22X1 U8928 ( .A0(n12398), .A1(n7940), .B0(test_se), .B1(n7380), .Y(n10121) );
  INVX1 U8929 ( .A(n10122), .Y(n6455) );
  AOI22X1 U8930 ( .A0(n12398), .A1(n8593), .B0(n12397), .B1(n7940), .Y(n10122)
         );
  INVX1 U8931 ( .A(n10123), .Y(n6454) );
  AOI22X1 U8932 ( .A0(n12397), .A1(n8593), .B0(n12399), .B1(n7940), .Y(n10123)
         );
  OAI21X1 U8933 ( .A0(n7869), .A1(n7751), .B0(n10124), .Y(n6453) );
  AOI22X1 U8934 ( .A0(n10125), .A1(n7940), .B0(n12383), .B1(n10126), .Y(n10124) );
  OAI21X1 U8935 ( .A0(test_se), .A1(n10127), .B0(n7919), .Y(n10126) );
  NOR2X1 U8936 ( .A(n12401), .B(n10128), .Y(n10125) );
  NAND3X1 U8937 ( .A(n10129), .B(n10130), .C(n10131), .Y(n6452) );
  NAND2X1 U8938 ( .A(test_se), .B(n7442), .Y(n10131) );
  NAND4X1 U8939 ( .A(n8357), .B(n7940), .C(n10128), .D(n10132), .Y(n10130) );
  NOR2X1 U8940 ( .A(n10133), .B(n10134), .Y(n10132) );
  MX2X1 U8941 ( .A(n9057), .B(n9059), .S0(n7658), .Y(n10134) );
  NOR2X1 U8942 ( .A(n7545), .B(n7295), .Y(n9059) );
  NOR2X1 U8943 ( .A(n7295), .B(n12381), .Y(n9057) );
  MX2X1 U8944 ( .A(n9046), .B(n9056), .S0(n7627), .Y(n10133) );
  NOR2X1 U8945 ( .A(n7545), .B(n12382), .Y(n9056) );
  NOR2X1 U8946 ( .A(n12381), .B(n12382), .Y(n9046) );
  INVX1 U8947 ( .A(n10127), .Y(n10128) );
  NAND2X1 U8948 ( .A(n10135), .B(n12383), .Y(n10129) );
  AOI21X1 U8949 ( .A0(n8357), .A1(n10127), .B0(n7951), .Y(n10135) );
  NAND2X1 U8950 ( .A(n8344), .B(n8632), .Y(n10127) );
  INVX1 U8951 ( .A(n9028), .Y(n8357) );
  NAND2X1 U8952 ( .A(n6763), .B(n10136), .Y(n9028) );
  NAND3X1 U8953 ( .A(n8631), .B(n7442), .C(n10137), .Y(n10136) );
  NOR2X1 U8954 ( .A(n7380), .B(n13003), .Y(n8631) );
  OAI21X1 U8955 ( .A0(n7869), .A1(n7801), .B0(n10138), .Y(n6451) );
  AOI21X1 U8956 ( .A0(n10117), .A1(n7246), .B0(n10139), .Y(n10138) );
  AOI21X1 U8957 ( .A0(n7921), .A1(n10140), .B0(n12997), .Y(n10139) );
  NAND3X1 U8958 ( .A(n10120), .B(n7869), .C(n10141), .Y(n10140) );
  OAI21X1 U8959 ( .A0(n13001), .A1(n7940), .B0(n10142), .Y(n6450) );
  MX2X1 U8960 ( .A(n10120), .B(n10143), .S0(n7249), .Y(n10142) );
  INVX1 U8961 ( .A(n10144), .Y(n6449) );
  AOI22X1 U8962 ( .A0(n10145), .A1(n10117), .B0(test_se), .B1(n7249), .Y(
        n10144) );
  XOR2X1 U8963 ( .A(n7354), .B(n9016), .Y(n10145) );
  OAI21X1 U8964 ( .A0(n13000), .A1(n7940), .B0(n10146), .Y(n6448) );
  MX2X1 U8965 ( .A(n10147), .B(n10148), .S0(n7255), .Y(n10146) );
  NAND2X1 U8966 ( .A(n10117), .B(n10149), .Y(n10148) );
  INVX1 U8967 ( .A(n10143), .Y(n10117) );
  NAND2X1 U8968 ( .A(n7940), .B(n10120), .Y(n10143) );
  NAND2X1 U8969 ( .A(n10141), .B(n10120), .Y(n10147) );
  NAND2X1 U8970 ( .A(n10141), .B(n7246), .Y(n10120) );
  INVX1 U8971 ( .A(n10149), .Y(n10141) );
  NAND2X1 U8972 ( .A(n9016), .B(n7354), .Y(n10149) );
  NOR2X1 U8973 ( .A(n9018), .B(n7546), .Y(n9016) );
  INVX1 U8974 ( .A(n9022), .Y(n9018) );
  NOR2X1 U8975 ( .A(n9014), .B(n12996), .Y(n9022) );
  NAND2X1 U8976 ( .A(n12999), .B(n7360), .Y(n9014) );
  NAND2X1 U8977 ( .A(n10150), .B(n10151), .Y(n6447) );
  AOI21X1 U8978 ( .A0(n10152), .A1(n8353), .B0(n10153), .Y(n10151) );
  AOI21X1 U8979 ( .A0(n10154), .A1(n10155), .B0(n12212), .Y(n10153) );
  NAND3X1 U8980 ( .A(n7940), .B(n10156), .C(n10157), .Y(n10155) );
  INVX1 U8981 ( .A(n8215), .Y(n10154) );
  INVX1 U8982 ( .A(n10157), .Y(n8353) );
  AOI21X1 U8983 ( .A0(n12327), .A1(n10158), .B0(n10159), .Y(n10157) );
  MX2X1 U8984 ( .A(n10160), .B(n10161), .S0(n7416), .Y(n10159) );
  NAND4X1 U8985 ( .A(n10162), .B(n10163), .C(n10164), .D(n10165), .Y(n10161)
         );
  NAND3X1 U8986 ( .A(n8220), .B(g17819), .C(n12323), .Y(n10165) );
  AOI22X1 U8987 ( .A0(n10166), .A1(n12325), .B0(n10167), .B1(n12324), .Y(
        n10164) );
  NOR2X1 U8988 ( .A(n5256), .B(n10168), .Y(n10167) );
  NOR2X1 U8989 ( .A(n7618), .B(n10169), .Y(n10166) );
  OR2X1 U8990 ( .A(n10170), .B(n10171), .Y(n10163) );
  AOI22X1 U8991 ( .A0(n12313), .A1(g13068), .B0(n12314), .B1(n12315), .Y(
        n10170) );
  MX2X1 U8992 ( .A(n10172), .B(n10173), .S0(g12350), .Y(n10162) );
  AOI21X1 U8993 ( .A0(n8220), .A1(n7443), .B0(n10174), .Y(n10173) );
  INVX1 U8994 ( .A(n10175), .Y(n10172) );
  NAND4X1 U8995 ( .A(n10176), .B(n10177), .C(n10178), .D(n10179), .Y(n10160)
         );
  OR2X1 U8996 ( .A(n10180), .B(n10168), .Y(n10179) );
  INVX1 U8997 ( .A(n8222), .Y(n10168) );
  AOI22X1 U8998 ( .A0(n12309), .A1(g13068), .B0(n12310), .B1(n12315), .Y(
        n10180) );
  AOI22X1 U8999 ( .A0(n10181), .A1(n12312), .B0(n10182), .B1(n12311), .Y(
        n10178) );
  NOR2X1 U9000 ( .A(n5257), .B(n10169), .Y(n10182) );
  INVX1 U9001 ( .A(n8221), .Y(n10169) );
  NOR2X1 U9002 ( .A(n5256), .B(n10171), .Y(n10181) );
  INVX1 U9003 ( .A(n8223), .Y(n10171) );
  OR2X1 U9004 ( .A(n10183), .B(n10184), .Y(n10177) );
  AOI22X1 U9005 ( .A0(n12308), .A1(g17715), .B0(n12307), .B1(g17646), .Y(
        n10183) );
  MX2X1 U9006 ( .A(n10185), .B(n10186), .S0(g12350), .Y(n10176) );
  AOI21X1 U9007 ( .A0(n8221), .A1(n7389), .B0(n10175), .Y(n10186) );
  NAND3X1 U9008 ( .A(n10187), .B(n10188), .C(n10189), .Y(n10175) );
  NAND3X1 U9009 ( .A(n8220), .B(g17739), .C(n12320), .Y(n10189) );
  NAND3X1 U9010 ( .A(n8223), .B(g14738), .C(n12322), .Y(n10188) );
  NAND3X1 U9011 ( .A(n8222), .B(g17607), .C(n12321), .Y(n10187) );
  INVX1 U9012 ( .A(n10174), .Y(n10185) );
  NAND3X1 U9013 ( .A(n10190), .B(n10191), .C(n10192), .Y(n10174) );
  NAND3X1 U9014 ( .A(n8222), .B(g14738), .C(n12318), .Y(n10192) );
  NAND3X1 U9015 ( .A(n8223), .B(g17607), .C(n12317), .Y(n10191) );
  NOR2X1 U9016 ( .A(n7253), .B(n12377), .Y(n8223) );
  NAND3X1 U9017 ( .A(n8221), .B(g17739), .C(n12319), .Y(n10190) );
  INVX1 U9018 ( .A(n10156), .Y(n10158) );
  INVX1 U9019 ( .A(n10193), .Y(n10152) );
  AOI21X1 U9020 ( .A0(n12212), .A1(n8352), .B0(n10194), .Y(n10193) );
  AOI22X1 U9021 ( .A0(n12213), .A1(n7893), .B0(n12215), .B1(test_se), .Y(
        n10150) );
  OAI21X1 U9022 ( .A0(n10195), .A1(n7569), .B0(n10196), .Y(n6446) );
  MX2X1 U9023 ( .A(n10197), .B(n7331), .S0(n7960), .Y(n10196) );
  NAND2X1 U9024 ( .A(n8540), .B(n7569), .Y(n10197) );
  OAI21X1 U9025 ( .A0(n12207), .A1(n10198), .B0(n10199), .Y(n6445) );
  OAI21X1 U9026 ( .A0(n8276), .A1(n8593), .B0(n12208), .Y(n10199) );
  OAI21X1 U9027 ( .A0(n12691), .A1(n10198), .B0(n10200), .Y(n6444) );
  MX2X1 U9028 ( .A(n10201), .B(n10202), .S0(n12207), .Y(n10200) );
  NAND2X1 U9029 ( .A(n10194), .B(n7569), .Y(n10202) );
  INVX1 U9030 ( .A(n10203), .Y(n10194) );
  AOI21X1 U9031 ( .A0(n12208), .A1(n8276), .B0(n8593), .Y(n10201) );
  OAI21X1 U9032 ( .A0(n12691), .A1(n7940), .B0(n10204), .Y(n6443) );
  MX2X1 U9033 ( .A(n10198), .B(n10203), .S0(n7584), .Y(n10204) );
  NAND2X1 U9034 ( .A(n8276), .B(n7940), .Y(n10203) );
  NOR2X1 U9035 ( .A(n10156), .B(n10205), .Y(n8276) );
  AOI21X1 U9036 ( .A0(n10156), .A1(n7941), .B0(n8215), .Y(n10198) );
  NAND3X1 U9037 ( .A(g17646), .B(n7416), .C(n8221), .Y(n10156) );
  NOR2X1 U9038 ( .A(n7547), .B(n12378), .Y(n8221) );
  MX2X1 U9039 ( .A(n12205), .B(n12206), .S0(n10195), .Y(n6442) );
  OAI21X1 U9040 ( .A0(n10195), .A1(n7641), .B0(n10206), .Y(n6441) );
  MX2X1 U9041 ( .A(n10207), .B(n10208), .S0(n12205), .Y(n10206) );
  AOI21X1 U9042 ( .A0(n12206), .A1(n8540), .B0(n8593), .Y(n10208) );
  NAND3X1 U9043 ( .A(n7941), .B(n7584), .C(n8540), .Y(n10207) );
  INVX1 U9044 ( .A(n8488), .Y(n10195) );
  INVX1 U9045 ( .A(n10209), .Y(n6440) );
  AOI22X1 U9046 ( .A0(n12204), .A1(n10210), .B0(n12209), .B1(test_se), .Y(
        n10209) );
  NAND2X1 U9047 ( .A(n10211), .B(n10212), .Y(n6439) );
  MX2X1 U9048 ( .A(n10213), .B(n12204), .S0(n7960), .Y(n10211) );
  INVX1 U9049 ( .A(n10214), .Y(n6438) );
  AOI22X1 U9050 ( .A0(n10215), .A1(n7261), .B0(n7946), .B1(n7429), .Y(n10214)
         );
  OAI21X1 U9051 ( .A0(n12211), .A1(n10216), .B0(n10217), .Y(n6437) );
  OAI21X1 U9052 ( .A0(n12211), .A1(n7983), .B0(n12210), .Y(n10217) );
  INVX1 U9053 ( .A(n10210), .Y(n10216) );
  NAND2X1 U9054 ( .A(n10218), .B(n10219), .Y(n6436) );
  MX2X1 U9055 ( .A(n10220), .B(n12211), .S0(n7960), .Y(n10219) );
  AOI21X1 U9056 ( .A0(n10210), .A1(n12214), .B0(n10221), .Y(n10218) );
  NOR2X1 U9057 ( .A(n7983), .B(n12210), .Y(n10210) );
  OAI21X1 U9058 ( .A0(n8534), .A1(n10222), .B0(n10223), .Y(n6435) );
  MX2X1 U9059 ( .A(n10224), .B(n7483), .S0(n7960), .Y(n10223) );
  NAND2X1 U9060 ( .A(n12313), .B(n10222), .Y(n10224) );
  OR2X1 U9061 ( .A(n10225), .B(n10226), .Y(n10222) );
  NAND2X1 U9062 ( .A(n10227), .B(n10228), .Y(n6434) );
  MX2X1 U9063 ( .A(n10229), .B(n8534), .S0(n10230), .Y(n10228) );
  NOR2X1 U9064 ( .A(n7261), .B(n10220), .Y(n10230) );
  NAND2X1 U9065 ( .A(n12310), .B(n7941), .Y(n10229) );
  AOI22X1 U9066 ( .A0(n12308), .A1(n7893), .B0(test_se), .B1(n7389), .Y(n10227) );
  NAND2X1 U9067 ( .A(n10231), .B(n10232), .Y(n6433) );
  MX2X1 U9068 ( .A(n10233), .B(n8534), .S0(n10234), .Y(n10232) );
  NOR2X1 U9069 ( .A(n10225), .B(n10212), .Y(n10234) );
  NAND2X1 U9070 ( .A(n12323), .B(n7941), .Y(n10233) );
  AOI22X1 U9071 ( .A0(n12313), .A1(n7893), .B0(n12310), .B1(test_se), .Y(
        n10231) );
  NAND2X1 U9072 ( .A(n10235), .B(n10236), .Y(n6432) );
  MX2X1 U9073 ( .A(n10237), .B(n8534), .S0(n10238), .Y(n10236) );
  NOR2X1 U9074 ( .A(n10213), .B(n10225), .Y(n10238) );
  NAND2X1 U9075 ( .A(n12324), .B(n7941), .Y(n10237) );
  AOI22X1 U9076 ( .A0(n12323), .A1(n7893), .B0(n12322), .B1(test_se), .Y(
        n10235) );
  NAND2X1 U9077 ( .A(n10239), .B(n10240), .Y(n6431) );
  MX2X1 U9078 ( .A(n10241), .B(n8534), .S0(n10242), .Y(n10240) );
  NOR2X1 U9079 ( .A(n10243), .B(n10225), .Y(n10242) );
  NAND2X1 U9080 ( .A(n12325), .B(n7941), .Y(n10241) );
  AOI22X1 U9081 ( .A0(n12324), .A1(n7892), .B0(n12320), .B1(test_se), .Y(
        n10239) );
  NAND2X1 U9082 ( .A(n10244), .B(n10245), .Y(n6430) );
  MX2X1 U9083 ( .A(n10246), .B(n8534), .S0(n10247), .Y(n10245) );
  NOR2X1 U9084 ( .A(n7261), .B(n10225), .Y(n10247) );
  NAND2X1 U9085 ( .A(n12211), .B(n7483), .Y(n10225) );
  NAND2X1 U9086 ( .A(n12314), .B(n7941), .Y(n10246) );
  AOI22X1 U9087 ( .A0(n12325), .A1(n7892), .B0(test_se), .B1(n7443), .Y(n10244) );
  NAND2X1 U9088 ( .A(n10248), .B(n10249), .Y(n6429) );
  AOI22X1 U9089 ( .A0(n10250), .A1(n7941), .B0(n10251), .B1(n10252), .Y(n10249) );
  AOI21X1 U9090 ( .A0(n10252), .A1(n10253), .B0(n12316), .Y(n10250) );
  INVX1 U9091 ( .A(n10226), .Y(n10252) );
  AOI22X1 U9092 ( .A0(n12314), .A1(n7892), .B0(n12313), .B1(test_se), .Y(
        n10248) );
  NAND2X1 U9093 ( .A(n10254), .B(n10255), .Y(n6428) );
  AOI22X1 U9094 ( .A0(n10256), .A1(n12318), .B0(n10251), .B1(n10257), .Y(
        n10255) );
  AOI21X1 U9095 ( .A0(n10257), .A1(n10253), .B0(n7983), .Y(n10256) );
  AOI22X1 U9096 ( .A0(n7892), .A1(n7443), .B0(n12323), .B1(test_se), .Y(n10254) );
  NAND2X1 U9097 ( .A(n10258), .B(n10259), .Y(n6427) );
  AOI22X1 U9098 ( .A0(n10260), .A1(n12319), .B0(n10251), .B1(n10261), .Y(
        n10259) );
  AOI21X1 U9099 ( .A0(n10253), .A1(n10261), .B0(n7983), .Y(n10260) );
  INVX1 U9100 ( .A(n10213), .Y(n10261) );
  AOI22X1 U9101 ( .A0(n12318), .A1(n7892), .B0(n12324), .B1(test_se), .Y(
        n10258) );
  NAND2X1 U9102 ( .A(n10262), .B(n10263), .Y(n6426) );
  AOI22X1 U9103 ( .A0(n10264), .A1(n12317), .B0(n10251), .B1(n10215), .Y(
        n10263) );
  AOI21X1 U9104 ( .A0(n10253), .A1(n10215), .B0(n7983), .Y(n10264) );
  AOI22X1 U9105 ( .A0(n12319), .A1(n7892), .B0(n12325), .B1(test_se), .Y(
        n10262) );
  NAND2X1 U9106 ( .A(n10265), .B(n10266), .Y(n6425) );
  AOI22X1 U9107 ( .A0(n10267), .A1(n12307), .B0(n10251), .B1(n12210), .Y(
        n10266) );
  AND2X1 U9108 ( .A(n10253), .B(n8893), .Y(n10251) );
  NOR2X1 U9109 ( .A(n10221), .B(n7983), .Y(n10267) );
  AND2X1 U9110 ( .A(n10253), .B(n12210), .Y(n10221) );
  NOR2X1 U9111 ( .A(n12214), .B(n12211), .Y(n10253) );
  AOI22X1 U9112 ( .A0(n12317), .A1(n7892), .B0(n12309), .B1(test_se), .Y(
        n10265) );
  NAND2X1 U9113 ( .A(n10268), .B(n10269), .Y(n6424) );
  MX2X1 U9114 ( .A(n10270), .B(n8534), .S0(n10271), .Y(n10269) );
  NOR2X1 U9115 ( .A(n10220), .B(n10226), .Y(n10271) );
  NAND2X1 U9116 ( .A(n12309), .B(n7941), .Y(n10270) );
  AOI22X1 U9117 ( .A0(n12307), .A1(n7892), .B0(n12314), .B1(test_se), .Y(
        n10268) );
  NAND2X1 U9118 ( .A(n10272), .B(n10273), .Y(n6423) );
  MX2X1 U9119 ( .A(n10274), .B(n8534), .S0(n10275), .Y(n10273) );
  NOR2X1 U9120 ( .A(n10220), .B(n10212), .Y(n10275) );
  NAND2X1 U9121 ( .A(n12311), .B(n7941), .Y(n10274) );
  AOI22X1 U9122 ( .A0(n12309), .A1(n7892), .B0(n12318), .B1(test_se), .Y(
        n10272) );
  NAND2X1 U9123 ( .A(n10276), .B(n10277), .Y(n6422) );
  MX2X1 U9124 ( .A(n10278), .B(n8534), .S0(n10279), .Y(n10277) );
  NOR2X1 U9125 ( .A(n10213), .B(n10220), .Y(n10279) );
  NAND2X1 U9126 ( .A(n12312), .B(n7941), .Y(n10278) );
  AOI22X1 U9127 ( .A0(n12311), .A1(n7892), .B0(n12319), .B1(test_se), .Y(
        n10276) );
  NAND2X1 U9128 ( .A(n10280), .B(n10281), .Y(n6421) );
  MX2X1 U9129 ( .A(n10282), .B(n8534), .S0(n10283), .Y(n10281) );
  NOR2X1 U9130 ( .A(n10284), .B(n10226), .Y(n10283) );
  NAND3X1 U9131 ( .A(n12204), .B(n7261), .C(n12203), .Y(n10226) );
  NAND2X1 U9132 ( .A(n7941), .B(n7389), .Y(n10282) );
  AOI22X1 U9133 ( .A0(n12310), .A1(n7892), .B0(n12307), .B1(test_se), .Y(
        n10280) );
  NAND2X1 U9134 ( .A(n10285), .B(n10286), .Y(n6420) );
  MX2X1 U9135 ( .A(n10287), .B(n8534), .S0(n10288), .Y(n10286) );
  NOR2X1 U9136 ( .A(n10284), .B(n10212), .Y(n10288) );
  INVX1 U9137 ( .A(n10257), .Y(n10212) );
  NOR2X1 U9138 ( .A(n7429), .B(n12204), .Y(n10257) );
  NAND2X1 U9139 ( .A(n12322), .B(n7941), .Y(n10287) );
  AOI22X1 U9140 ( .A0(n7892), .A1(n7389), .B0(n12311), .B1(test_se), .Y(n10285) );
  NAND2X1 U9141 ( .A(n10289), .B(n10290), .Y(n6419) );
  MX2X1 U9142 ( .A(n10291), .B(n8534), .S0(n10292), .Y(n10290) );
  NOR2X1 U9143 ( .A(n10284), .B(n10213), .Y(n10292) );
  NAND2X1 U9144 ( .A(n12204), .B(n7429), .Y(n10213) );
  NAND2X1 U9145 ( .A(n12320), .B(n7941), .Y(n10291) );
  AOI22X1 U9146 ( .A0(n12322), .A1(n7891), .B0(n12312), .B1(test_se), .Y(
        n10289) );
  NAND2X1 U9147 ( .A(n10293), .B(n10294), .Y(n6418) );
  MX2X1 U9148 ( .A(n10295), .B(n8534), .S0(n10296), .Y(n10294) );
  NOR2X1 U9149 ( .A(n10243), .B(n10220), .Y(n10296) );
  NAND2X1 U9150 ( .A(n12211), .B(n12214), .Y(n10220) );
  NAND2X1 U9151 ( .A(n12308), .B(n7941), .Y(n10295) );
  AOI22X1 U9152 ( .A0(n12312), .A1(n7891), .B0(n12317), .B1(test_se), .Y(
        n10293) );
  NAND2X1 U9153 ( .A(n10297), .B(n10298), .Y(n6417) );
  MX2X1 U9154 ( .A(n10299), .B(n8534), .S0(n10300), .Y(n10298) );
  NOR2X1 U9155 ( .A(n10284), .B(n10243), .Y(n10300) );
  INVX1 U9156 ( .A(n10215), .Y(n10243) );
  NOR2X1 U9157 ( .A(n12204), .B(n12203), .Y(n10215) );
  NAND2X1 U9158 ( .A(n12321), .B(n7941), .Y(n10299) );
  AOI22X1 U9159 ( .A0(n12320), .A1(n7891), .B0(n12308), .B1(test_se), .Y(
        n10297) );
  OAI21X1 U9160 ( .A0(n7941), .A1(n7802), .B0(n10301), .Y(n6416) );
  AOI22X1 U9161 ( .A0(n8488), .A1(n12327), .B0(n8893), .B1(n8540), .Y(n10301)
         );
  NOR2X1 U9162 ( .A(n7983), .B(n8540), .Y(n8488) );
  NOR2X1 U9163 ( .A(n7261), .B(n10284), .Y(n8540) );
  OR2X1 U9164 ( .A(n7483), .B(n12211), .Y(n10284) );
  MX2X1 U9165 ( .A(n12327), .B(g17739), .S0(n7848), .Y(n6415) );
  INVX1 U9166 ( .A(n10302), .Y(n6414) );
  MX2X1 U9167 ( .A(n10303), .B(n7869), .S0(g13068), .Y(n10302) );
  NAND4X1 U9168 ( .A(n7813), .B(n5568), .C(n10304), .D(n7941), .Y(n10303) );
  MX2X1 U9169 ( .A(n5569), .B(g12350), .S0(g14738), .Y(n10304) );
  MX2X1 U9170 ( .A(g17646), .B(g12350), .S0(n7848), .Y(n6413) );
  MX2X1 U9171 ( .A(g12350), .B(g14738), .S0(n7848), .Y(n6412) );
  OAI21X1 U9172 ( .A0(n10305), .A1(n10306), .B0(n10307), .Y(n6411) );
  MX2X1 U9173 ( .A(n10308), .B(n7803), .S0(n7960), .Y(n10307) );
  NAND2X1 U9174 ( .A(n10305), .B(n12326), .Y(n10308) );
  INVX1 U9175 ( .A(n10309), .Y(n10305) );
  OAI21X1 U9176 ( .A0(n7992), .A1(n7869), .B0(n10310), .Y(n6410) );
  AOI21X1 U9177 ( .A0(n12216), .A1(n7891), .B0(n10311), .Y(n10310) );
  INVX1 U9178 ( .A(n10312), .Y(n6409) );
  AOI22X1 U9179 ( .A0(n12214), .A1(n7941), .B0(n12216), .B1(test_se), .Y(
        n10312) );
  NOR2X1 U9180 ( .A(n10313), .B(n10314), .Y(n6408) );
  MX2X1 U9181 ( .A(n12376), .B(n12326), .S0(n7959), .Y(n10314) );
  NOR2X1 U9182 ( .A(n10313), .B(n7659), .Y(n6407) );
  NOR2X1 U9183 ( .A(n10306), .B(n10309), .Y(n10313) );
  NAND4X1 U9184 ( .A(g14738), .B(g17607), .C(g17739), .D(g12350), .Y(n10309)
         );
  INVX1 U9185 ( .A(n10311), .Y(n10306) );
  NOR2X1 U9186 ( .A(n7983), .B(n12326), .Y(n10311) );
  INVX1 U9187 ( .A(n10315), .Y(n6406) );
  AOI21X1 U9188 ( .A0(n7983), .A1(n12376), .B0(n10316), .Y(n10315) );
  MX2X1 U9189 ( .A(n8352), .B(n8215), .S0(n7253), .Y(n10316) );
  NOR2X1 U9190 ( .A(n10205), .B(n7983), .Y(n8352) );
  NAND2X1 U9191 ( .A(n10317), .B(n10318), .Y(n6405) );
  AOI22X1 U9192 ( .A0(n8222), .A1(n7941), .B0(n8215), .B1(n12377), .Y(n10318)
         );
  NOR2X1 U9193 ( .A(n7983), .B(n8219), .Y(n8215) );
  INVX1 U9194 ( .A(n10205), .Y(n8219) );
  NOR2X1 U9195 ( .A(n7547), .B(n7253), .Y(n8222) );
  AOI21X1 U9196 ( .A0(n7891), .A1(n7253), .B0(n10319), .Y(n10317) );
  MX2X1 U9197 ( .A(g14738), .B(n10320), .S0(n7848), .Y(n10319) );
  NOR2X1 U9198 ( .A(n10184), .B(n10205), .Y(n10320) );
  NAND2X1 U9199 ( .A(n4749), .B(n10321), .Y(n10205) );
  NAND3X1 U9200 ( .A(n12402), .B(n8345), .C(n10137), .Y(n10321) );
  NOR2X1 U9201 ( .A(n7249), .B(n13004), .Y(n8345) );
  INVX1 U9202 ( .A(n8220), .Y(n10184) );
  NOR2X1 U9203 ( .A(n12377), .B(n12378), .Y(n8220) );
  MX2X1 U9204 ( .A(n12377), .B(g17646), .S0(n7848), .Y(n6404) );
  NAND2X1 U9205 ( .A(n10322), .B(n10323), .Y(n6403) );
  AOI21X1 U9206 ( .A0(n10324), .A1(n9153), .B0(n10325), .Y(n10323) );
  AOI21X1 U9207 ( .A0(n8264), .A1(n10326), .B0(n12198), .Y(n10325) );
  NAND3X1 U9208 ( .A(n7941), .B(n10327), .C(n10328), .Y(n10326) );
  INVX1 U9209 ( .A(n10328), .Y(n9153) );
  AOI21X1 U9210 ( .A0(n12350), .A1(n10329), .B0(n10330), .Y(n10328) );
  MX2X1 U9211 ( .A(n10331), .B(n10332), .S0(n7417), .Y(n10330) );
  NAND4X1 U9212 ( .A(n10333), .B(n10334), .C(n10335), .D(n10336), .Y(n10332)
         );
  NAND3X1 U9213 ( .A(n10337), .B(g17845), .C(n12346), .Y(n10336) );
  AOI22X1 U9214 ( .A0(n10338), .A1(n12348), .B0(n10339), .B1(n12347), .Y(
        n10335) );
  NOR2X1 U9215 ( .A(n5254), .B(n8267), .Y(n10339) );
  NOR2X1 U9216 ( .A(n7596), .B(n8270), .Y(n10338) );
  OR2X1 U9217 ( .A(n10340), .B(n8268), .Y(n10334) );
  AOI22X1 U9218 ( .A0(n12336), .A1(g13085), .B0(n12337), .B1(n12338), .Y(
        n10340) );
  MX2X1 U9219 ( .A(n10341), .B(n10342), .S0(g12422), .Y(n10333) );
  AOI21X1 U9220 ( .A0(n10337), .A1(n7444), .B0(n10343), .Y(n10342) );
  INVX1 U9221 ( .A(n10344), .Y(n10341) );
  NAND4X1 U9222 ( .A(n10345), .B(n10346), .C(n10347), .D(n10348), .Y(n10331)
         );
  OR2X1 U9223 ( .A(n10349), .B(n8267), .Y(n10348) );
  INVX1 U9224 ( .A(n10350), .Y(n8267) );
  AOI22X1 U9225 ( .A0(n12332), .A1(g13085), .B0(n12333), .B1(n12338), .Y(
        n10349) );
  AOI22X1 U9226 ( .A0(n10351), .A1(n12335), .B0(n10352), .B1(n12334), .Y(
        n10347) );
  NOR2X1 U9227 ( .A(n5255), .B(n8270), .Y(n10352) );
  INVX1 U9228 ( .A(n10353), .Y(n8270) );
  NOR2X1 U9229 ( .A(n5254), .B(n8268), .Y(n10351) );
  INVX1 U9230 ( .A(n10354), .Y(n8268) );
  OR2X1 U9231 ( .A(n10355), .B(n8269), .Y(n10346) );
  AOI22X1 U9232 ( .A0(n12331), .A1(g17743), .B0(n12330), .B1(g17685), .Y(
        n10355) );
  MX2X1 U9233 ( .A(n10356), .B(n10357), .S0(g12422), .Y(n10345) );
  AOI21X1 U9234 ( .A0(n10353), .A1(n7390), .B0(n10344), .Y(n10357) );
  NAND3X1 U9235 ( .A(n10358), .B(n10359), .C(n10360), .Y(n10344) );
  NAND3X1 U9236 ( .A(n10337), .B(g17760), .C(n12343), .Y(n10360) );
  NAND3X1 U9237 ( .A(n10354), .B(g14779), .C(n12345), .Y(n10359) );
  NAND3X1 U9238 ( .A(n10350), .B(g17649), .C(n12344), .Y(n10358) );
  INVX1 U9239 ( .A(n10343), .Y(n10356) );
  NAND3X1 U9240 ( .A(n10361), .B(n10362), .C(n10363), .Y(n10343) );
  NAND3X1 U9241 ( .A(n10350), .B(g14779), .C(n12341), .Y(n10363) );
  NAND3X1 U9242 ( .A(n10354), .B(g17649), .C(n12340), .Y(n10362) );
  NOR2X1 U9243 ( .A(n7254), .B(n12373), .Y(n10354) );
  NAND3X1 U9244 ( .A(n10353), .B(g17760), .C(n12342), .Y(n10361) );
  INVX1 U9245 ( .A(n10327), .Y(n10329) );
  INVX1 U9246 ( .A(n10364), .Y(n10324) );
  AOI21X1 U9247 ( .A0(n8261), .A1(n12198), .B0(n10365), .Y(n10364) );
  AOI22X1 U9248 ( .A0(n12199), .A1(n7891), .B0(n12201), .B1(test_se), .Y(
        n10322) );
  OAI21X1 U9249 ( .A0(n10366), .A1(n7570), .B0(n10367), .Y(n6402) );
  MX2X1 U9250 ( .A(n10368), .B(n7621), .S0(n7959), .Y(n10367) );
  NAND2X1 U9251 ( .A(n8537), .B(n7570), .Y(n10368) );
  OAI21X1 U9252 ( .A0(n12193), .A1(n8306), .B0(n10369), .Y(n6401) );
  OAI21X1 U9253 ( .A0(n8311), .A1(n8593), .B0(n12194), .Y(n10369) );
  OAI21X1 U9254 ( .A0(n12690), .A1(n8306), .B0(n10370), .Y(n6400) );
  MX2X1 U9255 ( .A(n10371), .B(n10372), .S0(n12193), .Y(n10370) );
  NAND2X1 U9256 ( .A(n10365), .B(n7570), .Y(n10372) );
  INVX1 U9257 ( .A(n10373), .Y(n10365) );
  AOI21X1 U9258 ( .A0(n12194), .A1(n8311), .B0(n8593), .Y(n10371) );
  OAI21X1 U9259 ( .A0(n12690), .A1(n7941), .B0(n10374), .Y(n6399) );
  MX2X1 U9260 ( .A(n8306), .B(n10373), .S0(n7585), .Y(n10374) );
  NAND2X1 U9261 ( .A(n8311), .B(n7941), .Y(n10373) );
  OR2X1 U9262 ( .A(n7983), .B(n8311), .Y(n8306) );
  NOR2X1 U9263 ( .A(n10327), .B(n10375), .Y(n8311) );
  NAND3X1 U9264 ( .A(g17685), .B(n7417), .C(n10353), .Y(n10327) );
  NOR2X1 U9265 ( .A(n7548), .B(n12374), .Y(n10353) );
  MX2X1 U9266 ( .A(n12191), .B(n12192), .S0(n10366), .Y(n6398) );
  OAI21X1 U9267 ( .A0(n10366), .A1(n7642), .B0(n10376), .Y(n6397) );
  MX2X1 U9268 ( .A(n10377), .B(n10378), .S0(n12191), .Y(n10376) );
  AOI21X1 U9269 ( .A0(n12192), .A1(n8537), .B0(n8593), .Y(n10378) );
  NAND3X1 U9270 ( .A(n7941), .B(n7585), .C(n8537), .Y(n10377) );
  INVX1 U9271 ( .A(n8484), .Y(n10366) );
  INVX1 U9272 ( .A(n10379), .Y(n6396) );
  AOI22X1 U9273 ( .A0(n12190), .A1(n10380), .B0(n12195), .B1(test_se), .Y(
        n10379) );
  NAND2X1 U9274 ( .A(n10381), .B(n10382), .Y(n6395) );
  MX2X1 U9275 ( .A(n10383), .B(n12190), .S0(n7959), .Y(n10381) );
  INVX1 U9276 ( .A(n10384), .Y(n6394) );
  AOI22X1 U9277 ( .A0(n10385), .A1(n7262), .B0(n7983), .B1(n7430), .Y(n10384)
         );
  OAI21X1 U9278 ( .A0(n12197), .A1(n10386), .B0(n10387), .Y(n6393) );
  OAI21X1 U9279 ( .A0(n12197), .A1(n7982), .B0(n12196), .Y(n10387) );
  INVX1 U9280 ( .A(n10380), .Y(n10386) );
  NAND2X1 U9281 ( .A(n10388), .B(n10389), .Y(n6392) );
  MX2X1 U9282 ( .A(n10390), .B(n12197), .S0(n7957), .Y(n10389) );
  AOI21X1 U9283 ( .A0(n10380), .A1(n12200), .B0(n10391), .Y(n10388) );
  NOR2X1 U9284 ( .A(n7982), .B(n12196), .Y(n10380) );
  OAI21X1 U9285 ( .A0(n8534), .A1(n10392), .B0(n10393), .Y(n6391) );
  MX2X1 U9286 ( .A(n10394), .B(n7484), .S0(n7957), .Y(n10393) );
  NAND2X1 U9287 ( .A(n12336), .B(n10392), .Y(n10394) );
  OR2X1 U9288 ( .A(n10395), .B(n10396), .Y(n10392) );
  NAND2X1 U9289 ( .A(n10397), .B(n10398), .Y(n6390) );
  MX2X1 U9290 ( .A(n10399), .B(n8534), .S0(n10400), .Y(n10398) );
  NOR2X1 U9291 ( .A(n7262), .B(n10390), .Y(n10400) );
  NAND2X1 U9292 ( .A(n12333), .B(n7942), .Y(n10399) );
  AOI22X1 U9293 ( .A0(n12331), .A1(n7891), .B0(test_se), .B1(n7390), .Y(n10397) );
  NAND2X1 U9294 ( .A(n10401), .B(n10402), .Y(n6389) );
  MX2X1 U9295 ( .A(n10403), .B(n8534), .S0(n10404), .Y(n10402) );
  NOR2X1 U9296 ( .A(n10395), .B(n10382), .Y(n10404) );
  NAND2X1 U9297 ( .A(n12346), .B(n7942), .Y(n10403) );
  AOI22X1 U9298 ( .A0(n12336), .A1(n7891), .B0(n12333), .B1(test_se), .Y(
        n10401) );
  NAND2X1 U9299 ( .A(n10405), .B(n10406), .Y(n6388) );
  MX2X1 U9300 ( .A(n10407), .B(n8534), .S0(n10408), .Y(n10406) );
  NOR2X1 U9301 ( .A(n10383), .B(n10395), .Y(n10408) );
  NAND2X1 U9302 ( .A(n12347), .B(n7942), .Y(n10407) );
  AOI22X1 U9303 ( .A0(n12346), .A1(n7891), .B0(n12345), .B1(test_se), .Y(
        n10405) );
  NAND2X1 U9304 ( .A(n10409), .B(n10410), .Y(n6387) );
  MX2X1 U9305 ( .A(n10411), .B(n8534), .S0(n10412), .Y(n10410) );
  NOR2X1 U9306 ( .A(n10413), .B(n10395), .Y(n10412) );
  NAND2X1 U9307 ( .A(n12348), .B(n7942), .Y(n10411) );
  AOI22X1 U9308 ( .A0(n12347), .A1(n7891), .B0(n12343), .B1(test_se), .Y(
        n10409) );
  NAND2X1 U9309 ( .A(n10414), .B(n10415), .Y(n6386) );
  MX2X1 U9310 ( .A(n10416), .B(n8534), .S0(n10417), .Y(n10415) );
  NOR2X1 U9311 ( .A(n7262), .B(n10395), .Y(n10417) );
  NAND2X1 U9312 ( .A(n12197), .B(n7484), .Y(n10395) );
  NAND2X1 U9313 ( .A(n12337), .B(n7942), .Y(n10416) );
  AOI22X1 U9314 ( .A0(n12348), .A1(n7891), .B0(test_se), .B1(n7444), .Y(n10414) );
  NAND2X1 U9315 ( .A(n10418), .B(n10419), .Y(n6385) );
  AOI22X1 U9316 ( .A0(n10420), .A1(n7942), .B0(n10421), .B1(n10422), .Y(n10419) );
  AOI21X1 U9317 ( .A0(n10422), .A1(n10423), .B0(n12339), .Y(n10420) );
  INVX1 U9318 ( .A(n10396), .Y(n10422) );
  AOI22X1 U9319 ( .A0(n12337), .A1(n7891), .B0(n12336), .B1(test_se), .Y(
        n10418) );
  NAND2X1 U9320 ( .A(n10424), .B(n10425), .Y(n6384) );
  AOI22X1 U9321 ( .A0(n10426), .A1(n12341), .B0(n10421), .B1(n10427), .Y(
        n10425) );
  AOI21X1 U9322 ( .A0(n10427), .A1(n10423), .B0(n7982), .Y(n10426) );
  AOI22X1 U9323 ( .A0(n7890), .A1(n7444), .B0(n12346), .B1(test_se), .Y(n10424) );
  NAND2X1 U9324 ( .A(n10428), .B(n10429), .Y(n6383) );
  AOI22X1 U9325 ( .A0(n10430), .A1(n12342), .B0(n10421), .B1(n10431), .Y(
        n10429) );
  AOI21X1 U9326 ( .A0(n10423), .A1(n10431), .B0(n7982), .Y(n10430) );
  INVX1 U9327 ( .A(n10383), .Y(n10431) );
  AOI22X1 U9328 ( .A0(n12341), .A1(n7890), .B0(n12347), .B1(test_se), .Y(
        n10428) );
  NAND2X1 U9329 ( .A(n10432), .B(n10433), .Y(n6382) );
  AOI22X1 U9330 ( .A0(n10434), .A1(n12340), .B0(n10421), .B1(n10385), .Y(
        n10433) );
  AOI21X1 U9331 ( .A0(n10423), .A1(n10385), .B0(n7982), .Y(n10434) );
  AOI22X1 U9332 ( .A0(n12342), .A1(n7890), .B0(n12348), .B1(test_se), .Y(
        n10432) );
  NAND2X1 U9333 ( .A(n10435), .B(n10436), .Y(n6381) );
  AOI22X1 U9334 ( .A0(n10437), .A1(n12330), .B0(n10421), .B1(n12196), .Y(
        n10436) );
  AND2X1 U9335 ( .A(n10423), .B(n8893), .Y(n10421) );
  NOR2X1 U9336 ( .A(n10391), .B(n7982), .Y(n10437) );
  AND2X1 U9337 ( .A(n10423), .B(n12196), .Y(n10391) );
  NOR2X1 U9338 ( .A(n12200), .B(n12197), .Y(n10423) );
  AOI22X1 U9339 ( .A0(n12340), .A1(n7890), .B0(n12332), .B1(test_se), .Y(
        n10435) );
  NAND2X1 U9340 ( .A(n10438), .B(n10439), .Y(n6380) );
  MX2X1 U9341 ( .A(n10440), .B(n8534), .S0(n10441), .Y(n10439) );
  NOR2X1 U9342 ( .A(n10390), .B(n10396), .Y(n10441) );
  NAND2X1 U9343 ( .A(n12332), .B(n7942), .Y(n10440) );
  AOI22X1 U9344 ( .A0(n12330), .A1(n7890), .B0(n12337), .B1(test_se), .Y(
        n10438) );
  NAND2X1 U9345 ( .A(n10442), .B(n10443), .Y(n6379) );
  MX2X1 U9346 ( .A(n10444), .B(n8534), .S0(n10445), .Y(n10443) );
  NOR2X1 U9347 ( .A(n10390), .B(n10382), .Y(n10445) );
  NAND2X1 U9348 ( .A(n12334), .B(n7942), .Y(n10444) );
  AOI22X1 U9349 ( .A0(n12332), .A1(n7890), .B0(n12341), .B1(test_se), .Y(
        n10442) );
  NAND2X1 U9350 ( .A(n10446), .B(n10447), .Y(n6378) );
  MX2X1 U9351 ( .A(n10448), .B(n8534), .S0(n10449), .Y(n10447) );
  NOR2X1 U9352 ( .A(n10383), .B(n10390), .Y(n10449) );
  NAND2X1 U9353 ( .A(n12335), .B(n7942), .Y(n10448) );
  AOI22X1 U9354 ( .A0(n12334), .A1(n7890), .B0(n12342), .B1(test_se), .Y(
        n10446) );
  NAND2X1 U9355 ( .A(n10450), .B(n10451), .Y(n6377) );
  MX2X1 U9356 ( .A(n10452), .B(n8534), .S0(n10453), .Y(n10451) );
  NOR2X1 U9357 ( .A(n10454), .B(n10396), .Y(n10453) );
  NAND3X1 U9358 ( .A(n12190), .B(n7262), .C(n12189), .Y(n10396) );
  NAND2X1 U9359 ( .A(n7942), .B(n7390), .Y(n10452) );
  AOI22X1 U9360 ( .A0(n12333), .A1(n7890), .B0(n12330), .B1(test_se), .Y(
        n10450) );
  NAND2X1 U9361 ( .A(n10455), .B(n10456), .Y(n6376) );
  MX2X1 U9362 ( .A(n10457), .B(n8534), .S0(n10458), .Y(n10456) );
  NOR2X1 U9363 ( .A(n10454), .B(n10382), .Y(n10458) );
  INVX1 U9364 ( .A(n10427), .Y(n10382) );
  NOR2X1 U9365 ( .A(n7430), .B(n12190), .Y(n10427) );
  NAND2X1 U9366 ( .A(n12345), .B(n7942), .Y(n10457) );
  AOI22X1 U9367 ( .A0(n7890), .A1(n7390), .B0(n12334), .B1(test_se), .Y(n10455) );
  NAND2X1 U9368 ( .A(n10459), .B(n10460), .Y(n6375) );
  MX2X1 U9369 ( .A(n10461), .B(n8534), .S0(n10462), .Y(n10460) );
  NOR2X1 U9370 ( .A(n10454), .B(n10383), .Y(n10462) );
  NAND2X1 U9371 ( .A(n12190), .B(n7430), .Y(n10383) );
  NAND2X1 U9372 ( .A(n12343), .B(n7942), .Y(n10461) );
  AOI22X1 U9373 ( .A0(n12345), .A1(n7890), .B0(n12335), .B1(test_se), .Y(
        n10459) );
  NAND2X1 U9374 ( .A(n10463), .B(n10464), .Y(n6374) );
  MX2X1 U9375 ( .A(n10465), .B(n8534), .S0(n10466), .Y(n10464) );
  NOR2X1 U9376 ( .A(n10413), .B(n10390), .Y(n10466) );
  NAND2X1 U9377 ( .A(n12197), .B(n12200), .Y(n10390) );
  NAND2X1 U9378 ( .A(n12331), .B(n7942), .Y(n10465) );
  AOI22X1 U9379 ( .A0(n12335), .A1(n7890), .B0(n12340), .B1(test_se), .Y(
        n10463) );
  NAND2X1 U9380 ( .A(n10467), .B(n10468), .Y(n6373) );
  MX2X1 U9381 ( .A(n10469), .B(n8534), .S0(n10470), .Y(n10468) );
  NOR2X1 U9382 ( .A(n10454), .B(n10413), .Y(n10470) );
  INVX1 U9383 ( .A(n10385), .Y(n10413) );
  NOR2X1 U9384 ( .A(n12190), .B(n12189), .Y(n10385) );
  INVX1 U9385 ( .A(n8893), .Y(n8534) );
  NAND2X1 U9386 ( .A(n12344), .B(n7942), .Y(n10469) );
  AOI22X1 U9387 ( .A0(n12343), .A1(n7890), .B0(n12331), .B1(test_se), .Y(
        n10467) );
  OAI21X1 U9388 ( .A0(n7942), .A1(n7804), .B0(n10471), .Y(n6372) );
  AOI22X1 U9389 ( .A0(n8893), .A1(n8537), .B0(n12350), .B1(n8484), .Y(n10471)
         );
  NOR2X1 U9390 ( .A(n7982), .B(n8537), .Y(n8484) );
  NOR2X1 U9391 ( .A(n7262), .B(n10454), .Y(n8537) );
  OR2X1 U9392 ( .A(n7484), .B(n12197), .Y(n10454) );
  NOR2X1 U9393 ( .A(n7982), .B(n8557), .Y(n8893) );
  NOR2X1 U9394 ( .A(n7516), .B(n12593), .Y(n8557) );
  MX2X1 U9395 ( .A(n12350), .B(g17760), .S0(n7848), .Y(n6371) );
  INVX1 U9396 ( .A(n10472), .Y(n6370) );
  MX2X1 U9397 ( .A(n10473), .B(n7869), .S0(g13085), .Y(n10472) );
  NAND4X1 U9398 ( .A(n7809), .B(n5537), .C(n10474), .D(n7942), .Y(n10473) );
  MX2X1 U9399 ( .A(n5538), .B(g12422), .S0(g14779), .Y(n10474) );
  MX2X1 U9400 ( .A(g17685), .B(g12422), .S0(n7848), .Y(n6369) );
  MX2X1 U9401 ( .A(g12422), .B(g14779), .S0(n7847), .Y(n6368) );
  OAI21X1 U9402 ( .A0(n10475), .A1(n10476), .B0(n10477), .Y(n6367) );
  MX2X1 U9403 ( .A(n10478), .B(n7806), .S0(n7955), .Y(n10477) );
  NAND2X1 U9404 ( .A(n10475), .B(n12349), .Y(n10478) );
  INVX1 U9405 ( .A(n10479), .Y(n10475) );
  OAI21X1 U9406 ( .A0(n7994), .A1(n7869), .B0(n10480), .Y(n6366) );
  AOI21X1 U9407 ( .A0(n12202), .A1(n7889), .B0(n10481), .Y(n10480) );
  INVX1 U9408 ( .A(n10482), .Y(n6365) );
  AOI22X1 U9409 ( .A0(n12200), .A1(n7942), .B0(n12202), .B1(test_se), .Y(
        n10482) );
  NOR2X1 U9410 ( .A(n10483), .B(n10484), .Y(n6364) );
  MX2X1 U9411 ( .A(n12372), .B(n12349), .S0(n7948), .Y(n10484) );
  NOR2X1 U9412 ( .A(n10483), .B(n7660), .Y(n6363) );
  NOR2X1 U9413 ( .A(n10476), .B(n10479), .Y(n10483) );
  NAND4X1 U9414 ( .A(g14779), .B(g17649), .C(g17760), .D(g12422), .Y(n10479)
         );
  INVX1 U9415 ( .A(n10481), .Y(n10476) );
  NOR2X1 U9416 ( .A(n7982), .B(n12349), .Y(n10481) );
  INVX1 U9417 ( .A(n10485), .Y(n6362) );
  AOI21X1 U9418 ( .A0(n7982), .A1(n12372), .B0(n10486), .Y(n10485) );
  MX2X1 U9419 ( .A(n8261), .B(n9154), .S0(n7254), .Y(n10486) );
  NOR2X1 U9420 ( .A(n10375), .B(n7982), .Y(n8261) );
  NAND2X1 U9421 ( .A(n10487), .B(n10488), .Y(n6361) );
  AOI22X1 U9422 ( .A0(n9154), .A1(n12373), .B0(n10350), .B1(n7942), .Y(n10488)
         );
  NOR2X1 U9423 ( .A(n7548), .B(n7254), .Y(n10350) );
  INVX1 U9424 ( .A(n8264), .Y(n9154) );
  NAND2X1 U9425 ( .A(n7942), .B(n10375), .Y(n8264) );
  AOI21X1 U9426 ( .A0(n7889), .A1(n7254), .B0(n10489), .Y(n10487) );
  MX2X1 U9427 ( .A(g14779), .B(n10490), .S0(n7847), .Y(n10489) );
  NOR2X1 U9428 ( .A(n10375), .B(n8269), .Y(n10490) );
  INVX1 U9429 ( .A(n10337), .Y(n8269) );
  NOR2X1 U9430 ( .A(n12373), .B(n12374), .Y(n10337) );
  NAND2X1 U9431 ( .A(n7360), .B(n10491), .Y(n10375) );
  NAND3X1 U9432 ( .A(n12400), .B(n8636), .C(n10137), .Y(n10491) );
  MX2X1 U9433 ( .A(n12373), .B(g17685), .S0(n7847), .Y(n6360) );
  OAI21X1 U9434 ( .A0(n12405), .A1(n7869), .B0(n10492), .Y(n6359) );
  AOI22X1 U9435 ( .A0(n10493), .A1(n13002), .B0(n10494), .B1(n7459), .Y(n10492) );
  OAI21X1 U9436 ( .A0(test_se), .A1(n10109), .B0(n7919), .Y(n10494) );
  NOR2X1 U9437 ( .A(n10107), .B(n7982), .Y(n10493) );
  INVX1 U9438 ( .A(n10109), .Y(n10107) );
  NAND2X1 U9439 ( .A(n8344), .B(n8636), .Y(n10109) );
  NOR2X1 U9440 ( .A(n13004), .B(n13003), .Y(n8636) );
  INVX1 U9441 ( .A(n8584), .Y(n8344) );
  NAND3X1 U9442 ( .A(n7246), .B(n7354), .C(n12997), .Y(n8584) );
  MX2X1 U9443 ( .A(n12993), .B(g17577), .S0(n7847), .Y(n6358) );
  OAI21X1 U9444 ( .A0(n5533), .A1(n7869), .B0(n10495), .Y(n6357) );
  AOI21X1 U9445 ( .A0(n10496), .A1(g20557), .B0(n10497), .Y(n10495) );
  AOI21X1 U9446 ( .A0(n7921), .A1(n10498), .B0(n12260), .Y(n10497) );
  NAND4X1 U9447 ( .A(n5532), .B(n12261), .C(n7243), .D(n7869), .Y(n10498) );
  OR2X1 U9448 ( .A(n10499), .B(n9948), .Y(n10496) );
  NOR2X1 U9449 ( .A(n7243), .B(n7982), .Y(n9948) );
  AOI21X1 U9450 ( .A0(n12261), .A1(n7498), .B0(n7981), .Y(n10499) );
  OAI21X1 U9451 ( .A0(n7869), .A1(n7549), .B0(n10500), .Y(n6356) );
  AOI22X1 U9452 ( .A0(n13049), .A1(n7889), .B0(n7942), .B1(g29215), .Y(n10500)
         );
  MX2X1 U9453 ( .A(g8416), .B(g12919), .S0(n7847), .Y(n6355) );
  OAI21X1 U9454 ( .A0(n5529), .A1(n7942), .B0(n10501), .Y(n6354) );
  NAND2X1 U9455 ( .A(n10502), .B(n10503), .Y(n6353) );
  MX2X1 U9456 ( .A(n10501), .B(n10504), .S0(n7933), .Y(n10503) );
  NAND2X1 U9457 ( .A(n7942), .B(g10500), .Y(n10504) );
  INVX1 U9458 ( .A(n10505), .Y(n10501) );
  AOI22X1 U9459 ( .A0(n7889), .A1(n7500), .B0(test_se), .B1(g12919), .Y(n10502) );
  OAI21X1 U9460 ( .A0(n7869), .A1(n7517), .B0(n10506), .Y(n6352) );
  AOI21X1 U9461 ( .A0(n13062), .A1(n7889), .B0(n10505), .Y(n10506) );
  NOR2X1 U9462 ( .A(n7981), .B(n5888), .Y(n10505) );
  OAI21X1 U9463 ( .A0(n7869), .A1(n7371), .B0(n10507), .Y(n6351) );
  AOI22X1 U9464 ( .A0(n7942), .A1(n10508), .B0(n13070), .B1(n7889), .Y(n10507)
         );
  XOR2X1 U9465 ( .A(n10509), .B(n10510), .Y(n10508) );
  NAND3X1 U9466 ( .A(n5530), .B(n10511), .C(n768), .Y(n10510) );
  INVX1 U9467 ( .A(n10512), .Y(n10511) );
  NAND3X1 U9468 ( .A(n8132), .B(n10513), .C(n8131), .Y(n10509) );
  MX2X1 U9469 ( .A(n13062), .B(g7916), .S0(n7847), .Y(n6350) );
  MX2X1 U9470 ( .A(n13074), .B(g8416), .S0(n7847), .Y(n6349) );
  OAI21X1 U9471 ( .A0(n10514), .A1(n7472), .B0(n10515), .Y(n6348) );
  NAND3X1 U9472 ( .A(n7943), .B(n10516), .C(n13065), .Y(n10515) );
  OAI21X1 U9473 ( .A0(n13073), .A1(n10517), .B0(n10518), .Y(n10516) );
  AOI21X1 U9474 ( .A0(n10519), .A1(n10518), .B0(n7981), .Y(n10514) );
  NOR2X1 U9475 ( .A(n13065), .B(n10517), .Y(n10519) );
  INVX1 U9476 ( .A(n10520), .Y(n6347) );
  AOI22X1 U9477 ( .A0(n10521), .A1(n7943), .B0(n13065), .B1(n8593), .Y(n10520)
         );
  MX2X1 U9478 ( .A(n10522), .B(n13064), .S0(n8698), .Y(n10521) );
  NOR2X1 U9479 ( .A(n13064), .B(n7382), .Y(n10522) );
  OAI21X1 U9480 ( .A0(n10523), .A1(n7715), .B0(n10524), .Y(n6346) );
  NAND3X1 U9481 ( .A(n10525), .B(n7445), .C(n7943), .Y(n10524) );
  OAI21X1 U9482 ( .A0(n13064), .A1(n7382), .B0(n8131), .Y(n10525) );
  AOI21X1 U9483 ( .A0(n10526), .A1(n13069), .B0(n7981), .Y(n10523) );
  NOR2X1 U9484 ( .A(n8698), .B(n7382), .Y(n10526) );
  OAI21X1 U9485 ( .A0(n7869), .A1(n7476), .B0(n10527), .Y(n6345) );
  AOI22X1 U9486 ( .A0(n10528), .A1(n13071), .B0(n13068), .B1(n10529), .Y(
        n10527) );
  OAI21X1 U9487 ( .A0(test_se), .A1(n8698), .B0(n7919), .Y(n10529) );
  INVX1 U9488 ( .A(n8131), .Y(n8698) );
  NOR2X1 U9489 ( .A(n10530), .B(n10531), .Y(n8131) );
  AOI21X1 U9490 ( .A0(n8700), .A1(n10532), .B0(n7981), .Y(n10528) );
  OAI21X1 U9491 ( .A0(n13072), .A1(n7472), .B0(n8701), .Y(n10532) );
  NAND2X1 U9492 ( .A(n10533), .B(n10534), .Y(n6344) );
  MX2X1 U9493 ( .A(n10535), .B(n10536), .S0(n7418), .Y(n10534) );
  NAND2X1 U9494 ( .A(n7943), .B(n10537), .Y(n10536) );
  NAND2X1 U9495 ( .A(n10538), .B(n10539), .Y(n10535) );
  AOI22X1 U9496 ( .A0(n13076), .A1(n7889), .B0(n13071), .B1(test_se), .Y(
        n10533) );
  NAND2X1 U9497 ( .A(n10540), .B(n10541), .Y(n6343) );
  NAND3X1 U9498 ( .A(n10542), .B(n7571), .C(n10538), .Y(n10541) );
  MX2X1 U9499 ( .A(n10543), .B(n13072), .S0(n7952), .Y(n10540) );
  NAND2X1 U9500 ( .A(n13067), .B(n10544), .Y(n10543) );
  NAND2X1 U9501 ( .A(n10545), .B(n10546), .Y(n6342) );
  NAND3X1 U9502 ( .A(n10518), .B(n7472), .C(n10538), .Y(n10546) );
  MX2X1 U9503 ( .A(n10547), .B(n7571), .S0(n7952), .Y(n10545) );
  OR2X1 U9504 ( .A(n7472), .B(n10518), .Y(n10547) );
  AOI21X1 U9505 ( .A0(n7571), .A1(n10548), .B0(n10544), .Y(n10518) );
  INVX1 U9506 ( .A(n10542), .Y(n10544) );
  AOI21X1 U9507 ( .A0(n10548), .A1(n13072), .B0(n10537), .Y(n10542) );
  INVX1 U9508 ( .A(n10539), .Y(n10537) );
  AOI21X1 U9509 ( .A0(n7476), .A1(n10548), .B0(n10531), .Y(n10539) );
  INVX1 U9510 ( .A(n10517), .Y(n10548) );
  NAND2X1 U9511 ( .A(n10549), .B(n10550), .Y(n6341) );
  MX2X1 U9512 ( .A(n10551), .B(n10552), .S0(n7476), .Y(n10550) );
  NAND2X1 U9513 ( .A(n10538), .B(n8700), .Y(n10552) );
  NOR2X1 U9514 ( .A(n10517), .B(n7981), .Y(n10538) );
  NAND3X1 U9515 ( .A(n8701), .B(n7609), .C(n10553), .Y(n10517) );
  MX2X1 U9516 ( .A(n13071), .B(n8699), .S0(n10530), .Y(n10553) );
  NAND3X1 U9517 ( .A(n13073), .B(n7418), .C(n13071), .Y(n8699) );
  NAND2X1 U9518 ( .A(n10554), .B(n7445), .Y(n8701) );
  NAND2X1 U9519 ( .A(n10531), .B(n7943), .Y(n10551) );
  AOI22X1 U9520 ( .A0(n13071), .A1(n7889), .B0(n13070), .B1(test_se), .Y(
        n10549) );
  INVX1 U9521 ( .A(n10555), .Y(n6340) );
  AOI22X1 U9522 ( .A0(n10556), .A1(n7943), .B0(test_se), .B1(n7445), .Y(n10555) );
  NOR2X1 U9523 ( .A(n13074), .B(n10557), .Y(n10556) );
  AOI22X1 U9524 ( .A0(n8705), .A1(n10512), .B0(n13063), .B1(n10558), .Y(n10557) );
  NOR2X1 U9525 ( .A(n13063), .B(n5888), .Y(n8705) );
  OAI21X1 U9526 ( .A0(n7869), .A1(n7610), .B0(n10559), .Y(n6339) );
  MX2X1 U9527 ( .A(n10560), .B(n10561), .S0(n7517), .Y(n10559) );
  NAND3X1 U9528 ( .A(n13074), .B(n7943), .C(n10562), .Y(n10561) );
  INVX1 U9529 ( .A(n10563), .Y(n10562) );
  AOI21X1 U9530 ( .A0(n10563), .A1(n7869), .B0(n7889), .Y(n10560) );
  NAND3X1 U9531 ( .A(n10513), .B(n10554), .C(n8132), .Y(n10563) );
  XOR2X1 U9532 ( .A(n13062), .B(n13074), .Y(n10513) );
  OAI21X1 U9533 ( .A0(n766), .A1(n7868), .B0(n10564), .Y(n6338) );
  AOI22X1 U9534 ( .A0(n10565), .A1(n7266), .B0(n13063), .B1(n7889), .Y(n10564)
         );
  MX2X1 U9535 ( .A(n10566), .B(n10567), .S0(n7533), .Y(n10565) );
  AND2X1 U9536 ( .A(n7868), .B(n10568), .Y(n10567) );
  NOR2X1 U9537 ( .A(n10568), .B(n7981), .Y(n10566) );
  NOR2X1 U9538 ( .A(n10558), .B(n7610), .Y(n10568) );
  NAND2X1 U9539 ( .A(g12919), .B(n10512), .Y(n10558) );
  NAND3X1 U9540 ( .A(n763), .B(n7517), .C(n766), .Y(n10512) );
  NAND2X1 U9541 ( .A(n10569), .B(n10570), .Y(n6337) );
  AOI22X1 U9542 ( .A0(n13055), .A1(n10571), .B0(n13056), .B1(n8689), .Y(n10570) );
  AOI22X1 U9543 ( .A0(n13017), .A1(n7889), .B0(n13054), .B1(test_se), .Y(
        n10569) );
  OAI21X1 U9544 ( .A0(n8721), .A1(n7752), .B0(n10572), .Y(n6336) );
  AOI22X1 U9545 ( .A0(n10573), .A1(n10574), .B0(n10575), .B1(n13050), .Y(
        n10572) );
  AOI21X1 U9546 ( .A0(n10576), .A1(n13051), .B0(n7981), .Y(n10575) );
  INVX1 U9547 ( .A(n10577), .Y(n10574) );
  AND2X1 U9548 ( .A(n10578), .B(n8689), .Y(n10573) );
  NAND2X1 U9549 ( .A(n10579), .B(n10580), .Y(n6335) );
  INVX1 U9550 ( .A(n10581), .Y(n10580) );
  MX2X1 U9551 ( .A(n8689), .B(n10571), .S0(n13053), .Y(n10581) );
  AOI22X1 U9552 ( .A0(n10582), .A1(n7943), .B0(test_se), .B1(g7916), .Y(n10579) );
  INVX1 U9553 ( .A(n10583), .Y(n10582) );
  NAND2X1 U9554 ( .A(n10584), .B(n10585), .Y(n6334) );
  MX2X1 U9555 ( .A(n7635), .B(n10586), .S0(n7847), .Y(n10585) );
  MX2X1 U9556 ( .A(n8690), .B(n10587), .S0(g7916), .Y(n10586) );
  AOI21X1 U9557 ( .A0(n13053), .A1(n7889), .B0(n10588), .Y(n10584) );
  AOI21X1 U9558 ( .A0(n10589), .A1(n10583), .B0(n7981), .Y(n10588) );
  NAND2X1 U9559 ( .A(n10590), .B(n10591), .Y(n6333) );
  AOI22X1 U9560 ( .A0(n10571), .A1(n13056), .B0(n8689), .B1(n13070), .Y(n10591) );
  NOR2X1 U9561 ( .A(n7981), .B(n763), .Y(n8689) );
  NOR2X1 U9562 ( .A(g7916), .B(n7981), .Y(n10571) );
  AOI22X1 U9563 ( .A0(n13054), .A1(n7888), .B0(n13053), .B1(test_se), .Y(
        n10590) );
  OAI21X1 U9564 ( .A0(n8721), .A1(n7690), .B0(n10592), .Y(n6332) );
  NAND3X1 U9565 ( .A(n10593), .B(n10583), .C(n7943), .Y(n10592) );
  XOR2X1 U9566 ( .A(n7518), .B(n10594), .Y(n10593) );
  OAI21X1 U9567 ( .A0(n7868), .A1(n7533), .B0(n10595), .Y(n6331) );
  AOI22X1 U9568 ( .A0(n10596), .A1(n10583), .B0(n13052), .B1(n7888), .Y(n10595) );
  NAND3X1 U9569 ( .A(n10578), .B(g7916), .C(n10597), .Y(n10583) );
  AOI21X1 U9570 ( .A0(n13050), .A1(n10589), .B0(n10577), .Y(n10597) );
  NAND2X1 U9571 ( .A(n8132), .B(n8694), .Y(n10578) );
  NAND4X1 U9572 ( .A(n10530), .B(n8700), .C(n13076), .D(n10598), .Y(n8694) );
  AND2X1 U9573 ( .A(n13067), .B(n13065), .Y(n10598) );
  INVX1 U9574 ( .A(n10531), .Y(n8700) );
  NOR2X1 U9575 ( .A(n13074), .B(n13075), .Y(n10531) );
  INVX1 U9576 ( .A(n10554), .Y(n10530) );
  XOR2X1 U9577 ( .A(n7494), .B(n7266), .Y(n10554) );
  MX2X1 U9578 ( .A(n10599), .B(n10600), .S0(n7628), .Y(n10596) );
  AND2X1 U9579 ( .A(n7868), .B(n10576), .Y(n10600) );
  NOR2X1 U9580 ( .A(n10576), .B(n7981), .Y(n10599) );
  NOR2X1 U9581 ( .A(n7518), .B(n10594), .Y(n10576) );
  NAND3X1 U9582 ( .A(n10577), .B(g7916), .C(n8244), .Y(n10594) );
  NAND3X1 U9583 ( .A(n13070), .B(n7752), .C(n13056), .Y(n10577) );
  OAI21X1 U9584 ( .A0(n7868), .A1(n7518), .B0(n10601), .Y(n6330) );
  MX2X1 U9585 ( .A(n10602), .B(n10603), .S0(n13048), .Y(n10601) );
  AOI21X1 U9586 ( .A0(n7532), .A1(n7868), .B0(n7888), .Y(n10603) );
  NAND2X1 U9587 ( .A(n13047), .B(n7943), .Y(n10602) );
  OAI21X1 U9588 ( .A0(n7868), .A1(n7532), .B0(n10604), .Y(n6329) );
  AOI22X1 U9589 ( .A0(n10605), .A1(n13049), .B0(n13016), .B1(n10606), .Y(
        n10604) );
  OAI21X1 U9590 ( .A0(n13049), .A1(n8133), .B0(n7919), .Y(n10606) );
  AND2X1 U9591 ( .A(n8133), .B(n7943), .Y(n10605) );
  OAI21X1 U9592 ( .A0(n7868), .A1(n7537), .B0(n10607), .Y(n6328) );
  AOI22X1 U9593 ( .A0(n10608), .A1(n7943), .B0(n13046), .B1(n7888), .Y(n10607)
         );
  MX2X1 U9594 ( .A(n10609), .B(n13016), .S0(n8133), .Y(n10608) );
  NAND2X1 U9595 ( .A(n13046), .B(n10610), .Y(n8133) );
  NOR2X1 U9596 ( .A(n13016), .B(n13049), .Y(n10609) );
  NAND2X1 U9597 ( .A(n10611), .B(n10612), .Y(n6327) );
  MX2X1 U9598 ( .A(n7636), .B(n10613), .S0(n7846), .Y(n10612) );
  NAND2X1 U9599 ( .A(n10610), .B(n7549), .Y(n10613) );
  AOI22X1 U9600 ( .A0(n13047), .A1(n7888), .B0(n10614), .B1(n13046), .Y(n10611) );
  NOR2X1 U9601 ( .A(n10610), .B(n7981), .Y(n10614) );
  AND2X1 U9602 ( .A(n13047), .B(n13048), .Y(n10610) );
  NAND3X1 U9603 ( .A(n10615), .B(n10616), .C(n10617), .Y(n6326) );
  AOI22X1 U9604 ( .A0(n13045), .A1(n7888), .B0(n13048), .B1(test_se), .Y(
        n10617) );
  NAND3X1 U9605 ( .A(n7943), .B(n10618), .C(n13044), .Y(n10616) );
  NAND3X1 U9606 ( .A(n10619), .B(g13259), .C(n10620), .Y(n10618) );
  INVX1 U9607 ( .A(n10621), .Y(n10620) );
  NAND3X1 U9608 ( .A(n8243), .B(n10621), .C(n10619), .Y(n10615) );
  XOR2X1 U9609 ( .A(n8241), .B(n7356), .Y(n10621) );
  NAND2X1 U9610 ( .A(n10622), .B(n10623), .Y(n6325) );
  MX2X1 U9611 ( .A(n7716), .B(n10624), .S0(n7846), .Y(n10623) );
  AOI22X1 U9612 ( .A0(n13045), .A1(n8474), .B0(n13040), .B1(n7888), .Y(n10622)
         );
  OAI22X1 U9613 ( .A0(n7868), .A1(n7611), .B0(n10625), .B1(n7980), .Y(n6324)
         );
  AOI22X1 U9614 ( .A0(n13043), .A1(n10624), .B0(n8476), .B1(n7272), .Y(n10625)
         );
  NAND2X1 U9615 ( .A(n13040), .B(n8476), .Y(n10624) );
  MX2X1 U9616 ( .A(n13043), .B(n13040), .S0(n8474), .Y(n6323) );
  NOR2X1 U9617 ( .A(n7980), .B(n8476), .Y(n8474) );
  NOR2X1 U9618 ( .A(n10626), .B(n768), .Y(n8476) );
  NAND2X1 U9619 ( .A(n10627), .B(n10628), .Y(n6322) );
  MX2X1 U9620 ( .A(n10629), .B(n10630), .S0(n7367), .Y(n10628) );
  NAND2X1 U9621 ( .A(n7943), .B(n10630), .Y(n10629) );
  NAND4X1 U9622 ( .A(n8246), .B(n13045), .C(n13039), .D(n7371), .Y(n10630) );
  NOR2X1 U9623 ( .A(n10589), .B(n768), .Y(n8246) );
  INVX1 U9624 ( .A(n8244), .Y(n10589) );
  AOI22X1 U9625 ( .A0(n13039), .A1(n7888), .B0(n13045), .B1(test_se), .Y(
        n10627) );
  NAND3X1 U9626 ( .A(n10631), .B(n10632), .C(n10633), .Y(n6321) );
  AOI22X1 U9627 ( .A0(n13038), .A1(n7888), .B0(test_se), .B1(g13259), .Y(
        n10633) );
  NAND3X1 U9628 ( .A(n7943), .B(n10634), .C(n13037), .Y(n10632) );
  NAND3X1 U9629 ( .A(n8691), .B(g13259), .C(n10635), .Y(n10634) );
  INVX1 U9630 ( .A(n10636), .Y(n10635) );
  NAND3X1 U9631 ( .A(n8243), .B(n10636), .C(n8691), .Y(n10631) );
  XOR2X1 U9632 ( .A(n8241), .B(n7282), .Y(n10636) );
  INVX1 U9633 ( .A(n8239), .Y(n8241) );
  NOR2X1 U9634 ( .A(n10637), .B(n13042), .Y(n8239) );
  INVX1 U9635 ( .A(n10638), .Y(n8243) );
  NAND4X1 U9636 ( .A(n7943), .B(g13259), .C(n7272), .D(n7679), .Y(n10638) );
  OAI21X1 U9637 ( .A0(n7943), .A1(n7807), .B0(n10639), .Y(n6320) );
  MX2X1 U9638 ( .A(n8438), .B(n13036), .S0(n10640), .Y(n10639) );
  NOR2X1 U9639 ( .A(n10641), .B(n10642), .Y(n10640) );
  NAND2X1 U9640 ( .A(n13037), .B(n13045), .Y(n10642) );
  NAND3X1 U9641 ( .A(g13259), .B(n7371), .C(n8691), .Y(n10641) );
  NAND2X1 U9642 ( .A(n10643), .B(n10644), .Y(n6319) );
  MX2X1 U9643 ( .A(n10645), .B(n10646), .S0(n7356), .Y(n10644) );
  NAND3X1 U9644 ( .A(n7371), .B(n7868), .C(n10647), .Y(n10646) );
  INVX1 U9645 ( .A(n10648), .Y(n10647) );
  OAI21X1 U9646 ( .A0(n13040), .A1(n10648), .B0(n7922), .Y(n10645) );
  NAND4X1 U9647 ( .A(n13044), .B(n13045), .C(n10619), .D(g13259), .Y(n10648)
         );
  AOI22X1 U9648 ( .A0(n13044), .A1(n7888), .B0(n13036), .B1(test_se), .Y(
        n10643) );
  MX2X1 U9649 ( .A(n13039), .B(g19334), .S0(n7846), .Y(n6318) );
  OAI21X1 U9650 ( .A0(n12941), .A1(n7868), .B0(n10649), .Y(n6317) );
  AOI22X1 U9651 ( .A0(n12944), .A1(n7888), .B0(n12896), .B1(n7943), .Y(n10649)
         );
  MX2X1 U9652 ( .A(g8475), .B(g12923), .S0(n7846), .Y(n6316) );
  OAI21X1 U9653 ( .A0(n7943), .A1(n7474), .B0(n10650), .Y(n6315) );
  NAND2X1 U9654 ( .A(n10651), .B(n10652), .Y(n6314) );
  MX2X1 U9655 ( .A(n10650), .B(n10653), .S0(n699), .Y(n10652) );
  NAND2X1 U9656 ( .A(n7943), .B(g10527), .Y(n10653) );
  INVX1 U9657 ( .A(n10654), .Y(n10650) );
  AOI22X1 U9658 ( .A0(n12895), .A1(n7888), .B0(test_se), .B1(g12923), .Y(
        n10651) );
  MX2X1 U9659 ( .A(n12951), .B(g7946), .S0(n7846), .Y(n6313) );
  MX2X1 U9660 ( .A(n12964), .B(g8475), .S0(n7846), .Y(n6312) );
  OAI21X1 U9661 ( .A0(n7868), .A1(n7478), .B0(n10655), .Y(n6311) );
  AOI21X1 U9662 ( .A0(n12951), .A1(n7887), .B0(n10654), .Y(n10655) );
  NOR2X1 U9663 ( .A(n7980), .B(n5511), .Y(n10654) );
  OAI21X1 U9664 ( .A0(n7868), .A1(n7372), .B0(n10656), .Y(n6310) );
  AOI22X1 U9665 ( .A0(n7943), .A1(n10657), .B0(n12966), .B1(n7887), .Y(n10656)
         );
  XOR2X1 U9666 ( .A(n10658), .B(n10659), .Y(n10657) );
  NAND3X1 U9667 ( .A(n8126), .B(n10660), .C(n8125), .Y(n10659) );
  NAND4X1 U9668 ( .A(n721), .B(n719), .C(n10661), .D(n716), .Y(n10658) );
  NOR2X1 U9669 ( .A(n12963), .B(g8475), .Y(n10661) );
  NAND2X1 U9670 ( .A(n10662), .B(n10663), .Y(n6309) );
  AOI22X1 U9671 ( .A0(n12948), .A1(n10664), .B0(n12967), .B1(n10665), .Y(
        n10663) );
  AOI22X1 U9672 ( .A0(n12965), .A1(n7887), .B0(n12972), .B1(test_se), .Y(
        n10662) );
  OAI21X1 U9673 ( .A0(n8721), .A1(n7753), .B0(n10666), .Y(n6308) );
  AOI22X1 U9674 ( .A0(n10667), .A1(n10668), .B0(n10669), .B1(n12945), .Y(
        n10666) );
  AOI21X1 U9675 ( .A0(n10670), .A1(n12946), .B0(n7980), .Y(n10669) );
  INVX1 U9676 ( .A(n10671), .Y(n10668) );
  AND2X1 U9677 ( .A(n10672), .B(n10665), .Y(n10667) );
  OAI21X1 U9678 ( .A0(n8721), .A1(n7689), .B0(n10673), .Y(n6307) );
  NAND3X1 U9679 ( .A(n10674), .B(n10675), .C(n7943), .Y(n10673) );
  XOR2X1 U9680 ( .A(n7519), .B(n10676), .Y(n10674) );
  OAI21X1 U9681 ( .A0(n7868), .A1(n7519), .B0(n10677), .Y(n6306) );
  MX2X1 U9682 ( .A(n10678), .B(n10679), .S0(n7313), .Y(n10677) );
  NAND2X1 U9683 ( .A(n12942), .B(n7943), .Y(n10679) );
  AOI21X1 U9684 ( .A0(n7527), .A1(n7868), .B0(n7887), .Y(n10678) );
  OAI21X1 U9685 ( .A0(n7868), .A1(n7527), .B0(n10680), .Y(n6305) );
  AOI22X1 U9686 ( .A0(n10681), .A1(n12944), .B0(n12897), .B1(n10682), .Y(
        n10680) );
  OAI21X1 U9687 ( .A0(n12944), .A1(n8127), .B0(n7919), .Y(n10682) );
  AND2X1 U9688 ( .A(n8127), .B(n7943), .Y(n10681) );
  OAI21X1 U9689 ( .A0(n7868), .A1(n7509), .B0(n10683), .Y(n6304) );
  AOI22X1 U9690 ( .A0(n10684), .A1(n7944), .B0(n7887), .B1(n7496), .Y(n10683)
         );
  MX2X1 U9691 ( .A(n10685), .B(n12897), .S0(n8127), .Y(n10684) );
  NAND2X1 U9692 ( .A(n10686), .B(n7496), .Y(n8127) );
  NOR2X1 U9693 ( .A(n12897), .B(n12944), .Y(n10685) );
  NAND2X1 U9694 ( .A(n10687), .B(n10688), .Y(n6303) );
  MX2X1 U9695 ( .A(n7637), .B(n10689), .S0(n7846), .Y(n10688) );
  NAND2X1 U9696 ( .A(n12941), .B(n10686), .Y(n10689) );
  AOI22X1 U9697 ( .A0(n12942), .A1(n7887), .B0(n10690), .B1(n7944), .Y(n10687)
         );
  NOR2X1 U9698 ( .A(n12941), .B(n10686), .Y(n10690) );
  NOR2X1 U9699 ( .A(n7527), .B(n7313), .Y(n10686) );
  NAND3X1 U9700 ( .A(n10691), .B(n10692), .C(n10693), .Y(n6302) );
  AOI22X1 U9701 ( .A0(n12971), .A1(n7887), .B0(n12943), .B1(test_se), .Y(
        n10693) );
  NAND4X1 U9702 ( .A(n10694), .B(n8232), .C(n10695), .D(g13272), .Y(n10692) );
  NAND3X1 U9703 ( .A(n7944), .B(n10696), .C(n12912), .Y(n10691) );
  NAND3X1 U9704 ( .A(n10694), .B(g13272), .C(n10697), .Y(n10696) );
  INVX1 U9705 ( .A(n10695), .Y(n10697) );
  XOR2X1 U9706 ( .A(n8230), .B(n12913), .Y(n10695) );
  NAND2X1 U9707 ( .A(n10698), .B(n10699), .Y(n6301) );
  INVX1 U9708 ( .A(n10700), .Y(n10699) );
  MX2X1 U9709 ( .A(n12912), .B(n10701), .S0(n7845), .Y(n10700) );
  AOI22X1 U9710 ( .A0(n10702), .A1(n12971), .B0(n12969), .B1(n7887), .Y(n10698) );
  OAI21X1 U9711 ( .A0(n7868), .A1(n7717), .B0(n10703), .Y(n6300) );
  AOI22X1 U9712 ( .A0(n10704), .A1(n12911), .B0(n8466), .B1(n10705), .Y(n10703) );
  NOR2X1 U9713 ( .A(n10701), .B(n7980), .Y(n10704) );
  AND2X1 U9714 ( .A(n12969), .B(n8466), .Y(n10701) );
  MX2X1 U9715 ( .A(n12911), .B(n12969), .S0(n10702), .Y(n6299) );
  NOR2X1 U9716 ( .A(n8466), .B(n7980), .Y(n10702) );
  NAND2X1 U9717 ( .A(n10706), .B(n10707), .Y(n6298) );
  MX2X1 U9718 ( .A(n13006), .B(n10708), .S0(n7845), .Y(n10707) );
  NAND3X1 U9719 ( .A(n12971), .B(n7534), .C(n10709), .Y(n10708) );
  AOI22X1 U9720 ( .A0(n12970), .A1(n7887), .B0(n12968), .B1(n10710), .Y(n10706) );
  OAI21X1 U9721 ( .A0(n10709), .A1(n7980), .B0(n10711), .Y(n10710) );
  INVX1 U9722 ( .A(n10712), .Y(n10709) );
  NAND3X1 U9723 ( .A(n8466), .B(n7372), .C(n12970), .Y(n10712) );
  AND2X1 U9724 ( .A(n10713), .B(g13272), .Y(n8466) );
  NAND2X1 U9725 ( .A(n10714), .B(n10715), .Y(n6297) );
  AOI22X1 U9726 ( .A0(n10716), .A1(n12965), .B0(n10717), .B1(n10665), .Y(
        n10715) );
  NOR2X1 U9727 ( .A(n7495), .B(n10718), .Y(n10717) );
  AOI21X1 U9728 ( .A0(n10719), .A1(g7946), .B0(n7980), .Y(n10716) );
  AOI22X1 U9729 ( .A0(n12967), .A1(n7887), .B0(n12968), .B1(test_se), .Y(
        n10714) );
  INVX1 U9730 ( .A(n10720), .Y(n6296) );
  AOI22X1 U9731 ( .A0(n7944), .A1(n10721), .B0(n12965), .B1(test_se), .Y(
        n10720) );
  OAI21X1 U9732 ( .A0(n12956), .A1(n10722), .B0(n10723), .Y(n10721) );
  AOI22X1 U9733 ( .A0(n10724), .A1(n10725), .B0(n12955), .B1(n10726), .Y(
        n10723) );
  INVX1 U9734 ( .A(n10727), .Y(n10725) );
  AND2X1 U9735 ( .A(n10728), .B(n10729), .Y(n10724) );
  OAI21X1 U9736 ( .A0(n7868), .A1(n7612), .B0(n10730), .Y(n6295) );
  AOI22X1 U9737 ( .A0(n7944), .A1(n10731), .B0(n12954), .B1(n10732), .Y(n10730) );
  OAI21X1 U9738 ( .A0(test_se), .A1(n5511), .B0(n7919), .Y(n10732) );
  OR2X1 U9739 ( .A(n10733), .B(n719), .Y(n10731) );
  AOI21X1 U9740 ( .A0(n7423), .A1(g12923), .B0(n12954), .Y(n10733) );
  MX2X1 U9741 ( .A(n12952), .B(g13272), .S0(n7845), .Y(n6294) );
  OAI21X1 U9742 ( .A0(n10734), .A1(n7473), .B0(n10735), .Y(n6293) );
  NAND3X1 U9743 ( .A(n7944), .B(n10736), .C(n12961), .Y(n10735) );
  OAI21X1 U9744 ( .A0(n12959), .A1(n10737), .B0(n10738), .Y(n10736) );
  AOI21X1 U9745 ( .A0(n10739), .A1(n10738), .B0(n7980), .Y(n10734) );
  NOR2X1 U9746 ( .A(n12961), .B(n10737), .Y(n10739) );
  INVX1 U9747 ( .A(n10740), .Y(n6292) );
  AOI22X1 U9748 ( .A0(n10741), .A1(n7944), .B0(n12961), .B1(n8593), .Y(n10740)
         );
  MX2X1 U9749 ( .A(n10742), .B(n12949), .S0(n10726), .Y(n10741) );
  NOR2X1 U9750 ( .A(n12949), .B(n7383), .Y(n10742) );
  OAI21X1 U9751 ( .A0(n10743), .A1(n7718), .B0(n10744), .Y(n6291) );
  NAND3X1 U9752 ( .A(n10745), .B(n7501), .C(n7944), .Y(n10744) );
  OAI21X1 U9753 ( .A0(n12949), .A1(n7383), .B0(n8125), .Y(n10745) );
  AOI21X1 U9754 ( .A0(n10746), .A1(n12957), .B0(n7980), .Y(n10743) );
  NOR2X1 U9755 ( .A(n10726), .B(n7383), .Y(n10746) );
  OAI21X1 U9756 ( .A0(n7868), .A1(n7477), .B0(n10747), .Y(n6290) );
  AOI22X1 U9757 ( .A0(n10748), .A1(n12956), .B0(n12955), .B1(n10749), .Y(
        n10747) );
  OAI21X1 U9758 ( .A0(test_se), .A1(n10726), .B0(n7919), .Y(n10749) );
  INVX1 U9759 ( .A(n8125), .Y(n10726) );
  NOR2X1 U9760 ( .A(n10750), .B(n10751), .Y(n8125) );
  AOI21X1 U9761 ( .A0(n10728), .A1(n10752), .B0(n7980), .Y(n10748) );
  OAI21X1 U9762 ( .A0(n12958), .A1(n7473), .B0(n10729), .Y(n10752) );
  NAND2X1 U9763 ( .A(n10753), .B(n10754), .Y(n6289) );
  MX2X1 U9764 ( .A(n10755), .B(n10756), .S0(n7477), .Y(n10754) );
  NAND2X1 U9765 ( .A(n10757), .B(n10728), .Y(n10756) );
  NAND2X1 U9766 ( .A(n10751), .B(n7944), .Y(n10755) );
  AOI22X1 U9767 ( .A0(n12956), .A1(n7887), .B0(n12966), .B1(test_se), .Y(
        n10753) );
  NAND2X1 U9768 ( .A(n10758), .B(n10759), .Y(n6288) );
  MX2X1 U9769 ( .A(n10760), .B(n10761), .S0(n7419), .Y(n10759) );
  NAND2X1 U9770 ( .A(n7944), .B(n10762), .Y(n10761) );
  NAND2X1 U9771 ( .A(n10757), .B(n10763), .Y(n10760) );
  AOI22X1 U9772 ( .A0(n12962), .A1(n7887), .B0(n12956), .B1(test_se), .Y(
        n10758) );
  NAND2X1 U9773 ( .A(n10764), .B(n10765), .Y(n6287) );
  NAND3X1 U9774 ( .A(n10766), .B(n7572), .C(n10757), .Y(n10765) );
  MX2X1 U9775 ( .A(n10767), .B(n12958), .S0(n7946), .Y(n10764) );
  NAND2X1 U9776 ( .A(n12960), .B(n10768), .Y(n10767) );
  NAND2X1 U9777 ( .A(n10769), .B(n10770), .Y(n6286) );
  NAND3X1 U9778 ( .A(n10738), .B(n7473), .C(n10757), .Y(n10770) );
  NOR2X1 U9779 ( .A(n10737), .B(n7980), .Y(n10757) );
  MX2X1 U9780 ( .A(n10771), .B(n7572), .S0(n7946), .Y(n10769) );
  OR2X1 U9781 ( .A(n7473), .B(n10738), .Y(n10771) );
  AOI21X1 U9782 ( .A0(n7572), .A1(n10772), .B0(n10768), .Y(n10738) );
  INVX1 U9783 ( .A(n10766), .Y(n10768) );
  AOI21X1 U9784 ( .A0(n10772), .A1(n12958), .B0(n10762), .Y(n10766) );
  INVX1 U9785 ( .A(n10763), .Y(n10762) );
  AOI21X1 U9786 ( .A0(n7477), .A1(n10772), .B0(n10751), .Y(n10763) );
  INVX1 U9787 ( .A(n10737), .Y(n10772) );
  NAND3X1 U9788 ( .A(n10729), .B(n7612), .C(n10773), .Y(n10737) );
  MX2X1 U9789 ( .A(n12956), .B(n10727), .S0(n10750), .Y(n10773) );
  NAND3X1 U9790 ( .A(n12959), .B(n7419), .C(n12956), .Y(n10727) );
  NAND2X1 U9791 ( .A(n10774), .B(n7501), .Y(n10729) );
  NAND2X1 U9792 ( .A(n10775), .B(n10776), .Y(n6285) );
  INVX1 U9793 ( .A(n10777), .Y(n10776) );
  MX2X1 U9794 ( .A(n10665), .B(n10664), .S0(n12973), .Y(n10777) );
  AOI22X1 U9795 ( .A0(n10778), .A1(n7944), .B0(test_se), .B1(g7946), .Y(n10775) );
  INVX1 U9796 ( .A(n10675), .Y(n10778) );
  NAND2X1 U9797 ( .A(n10779), .B(n10780), .Y(n6284) );
  MX2X1 U9798 ( .A(n7638), .B(n10781), .S0(n7845), .Y(n10780) );
  MX2X1 U9799 ( .A(n10718), .B(n10782), .S0(g7946), .Y(n10781) );
  AOI21X1 U9800 ( .A0(n12973), .A1(n7886), .B0(n10783), .Y(n10779) );
  AOI21X1 U9801 ( .A0(n10784), .A1(n10675), .B0(n7980), .Y(n10783) );
  NAND2X1 U9802 ( .A(n10785), .B(n10786), .Y(n6283) );
  AOI22X1 U9803 ( .A0(n12967), .A1(n10664), .B0(n10665), .B1(n12966), .Y(
        n10786) );
  NOR2X1 U9804 ( .A(n7979), .B(n716), .Y(n10665) );
  NOR2X1 U9805 ( .A(g7946), .B(n7979), .Y(n10664) );
  AOI22X1 U9806 ( .A0(n12972), .A1(n7886), .B0(n12973), .B1(test_se), .Y(
        n10785) );
  OAI21X1 U9807 ( .A0(n12957), .A1(n7868), .B0(n10787), .Y(n6282) );
  NAND3X1 U9808 ( .A(n10788), .B(n7256), .C(n7944), .Y(n10787) );
  XOR2X1 U9809 ( .A(n7423), .B(n10789), .Y(n10788) );
  OAI21X1 U9810 ( .A0(n7868), .A1(n7423), .B0(n10790), .Y(n6281) );
  MX2X1 U9811 ( .A(n10791), .B(n10792), .S0(n7478), .Y(n10790) );
  NAND3X1 U9812 ( .A(n12964), .B(n7944), .C(n10793), .Y(n10792) );
  INVX1 U9813 ( .A(n10794), .Y(n10793) );
  AOI21X1 U9814 ( .A0(n10794), .A1(n7868), .B0(n7886), .Y(n10791) );
  NAND3X1 U9815 ( .A(n10660), .B(n10774), .C(n8126), .Y(n10794) );
  XOR2X1 U9816 ( .A(n12951), .B(n12964), .Y(n10660) );
  MX2X1 U9817 ( .A(n12910), .B(g19357), .S0(n7845), .Y(n6280) );
  NAND2X1 U9818 ( .A(n10795), .B(n10796), .Y(n6279) );
  AOI22X1 U9819 ( .A0(n10797), .A1(n10798), .B0(n10799), .B1(n12907), .Y(
        n10796) );
  AOI21X1 U9820 ( .A0(n10800), .A1(n10798), .B0(n7979), .Y(n10799) );
  NOR2X1 U9821 ( .A(n10800), .B(n8469), .Y(n10797) );
  INVX1 U9822 ( .A(n8232), .Y(n8469) );
  NOR2X1 U9823 ( .A(n10711), .B(n12911), .Y(n8232) );
  INVX1 U9824 ( .A(n10705), .Y(n10711) );
  NOR2X1 U9825 ( .A(n7979), .B(n12971), .Y(n10705) );
  XOR2X1 U9826 ( .A(n8229), .B(n12908), .Y(n10800) );
  INVX1 U9827 ( .A(n8230), .Y(n8229) );
  NOR2X1 U9828 ( .A(n10801), .B(n12952), .Y(n8230) );
  AOI22X1 U9829 ( .A0(n12909), .A1(n7886), .B0(test_se), .B1(g13272), .Y(
        n10795) );
  OAI21X1 U9830 ( .A0(n12908), .A1(n10802), .B0(n10803), .Y(n6278) );
  MX2X1 U9831 ( .A(n10804), .B(n7808), .S0(n7953), .Y(n10803) );
  NAND2X1 U9832 ( .A(n12908), .B(n10802), .Y(n10804) );
  NAND4X1 U9833 ( .A(n12907), .B(n10798), .C(n12971), .D(n7372), .Y(n10802) );
  NOR2X1 U9834 ( .A(n10718), .B(n721), .Y(n10798) );
  NAND2X1 U9835 ( .A(n10805), .B(n10806), .Y(n6277) );
  MX2X1 U9836 ( .A(n10807), .B(n10808), .S0(n12913), .Y(n10806) );
  OAI21X1 U9837 ( .A0(n12969), .A1(n10809), .B0(n7923), .Y(n10808) );
  NAND3X1 U9838 ( .A(n7372), .B(n7868), .C(n10810), .Y(n10807) );
  INVX1 U9839 ( .A(n10809), .Y(n10810) );
  NAND4X1 U9840 ( .A(n12971), .B(n12912), .C(n10694), .D(g13272), .Y(n10809)
         );
  AOI22X1 U9841 ( .A0(n12912), .A1(n7886), .B0(n12908), .B1(test_se), .Y(
        n10805) );
  NAND2X1 U9842 ( .A(n10811), .B(n10812), .Y(n6276) );
  MX2X1 U9843 ( .A(n10813), .B(n10814), .S0(n12909), .Y(n10812) );
  NAND2X1 U9844 ( .A(n7944), .B(n10813), .Y(n10814) );
  NAND4X1 U9845 ( .A(n12971), .B(n8233), .C(n12910), .D(n7372), .Y(n10813) );
  NOR2X1 U9846 ( .A(n10784), .B(n721), .Y(n8233) );
  AOI22X1 U9847 ( .A0(n12910), .A1(n7886), .B0(n12971), .B1(test_se), .Y(
        n10811) );
  OAI21X1 U9848 ( .A0(n719), .A1(n7867), .B0(n10815), .Y(n6275) );
  AOI22X1 U9849 ( .A0(n10816), .A1(n7256), .B0(n12953), .B1(n7886), .Y(n10815)
         );
  MX2X1 U9850 ( .A(n10817), .B(n10818), .S0(n7479), .Y(n10816) );
  AND2X1 U9851 ( .A(n7867), .B(n10819), .Y(n10818) );
  NOR2X1 U9852 ( .A(n10819), .B(n7979), .Y(n10817) );
  NOR2X1 U9853 ( .A(n10789), .B(n7423), .Y(n10819) );
  NAND2X1 U9854 ( .A(g12923), .B(n10820), .Y(n10789) );
  NAND3X1 U9855 ( .A(n716), .B(n7478), .C(n719), .Y(n10820) );
  OAI21X1 U9856 ( .A0(n7867), .A1(n7479), .B0(n10821), .Y(n6274) );
  AOI22X1 U9857 ( .A0(n10822), .A1(n10675), .B0(n12947), .B1(n7886), .Y(n10821) );
  NAND3X1 U9858 ( .A(n10672), .B(g7946), .C(n10823), .Y(n10675) );
  AOI21X1 U9859 ( .A0(n12945), .A1(n10784), .B0(n10671), .Y(n10823) );
  INVX1 U9860 ( .A(n10824), .Y(n10784) );
  NAND2X1 U9861 ( .A(n8126), .B(n10722), .Y(n10672) );
  NAND4X1 U9862 ( .A(n10750), .B(n10728), .C(n12962), .D(n10825), .Y(n10722)
         );
  AND2X1 U9863 ( .A(n12961), .B(n12960), .Y(n10825) );
  INVX1 U9864 ( .A(n10751), .Y(n10728) );
  NOR2X1 U9865 ( .A(n12963), .B(n12964), .Y(n10751) );
  INVX1 U9866 ( .A(n10774), .Y(n10750) );
  XOR2X1 U9867 ( .A(n7495), .B(n7256), .Y(n10774) );
  MX2X1 U9868 ( .A(n10826), .B(n10827), .S0(n7629), .Y(n10822) );
  AND2X1 U9869 ( .A(n7867), .B(n10670), .Y(n10827) );
  NOR2X1 U9870 ( .A(n10670), .B(n7979), .Y(n10826) );
  NOR2X1 U9871 ( .A(n7519), .B(n10676), .Y(n10670) );
  NAND3X1 U9872 ( .A(n10671), .B(g7946), .C(n10824), .Y(n10676) );
  NAND3X1 U9873 ( .A(n12966), .B(n7753), .C(n12967), .Y(n10671) );
  NAND2X1 U9874 ( .A(n10828), .B(n10829), .Y(n6273) );
  AOI22X1 U9875 ( .A0(n12926), .A1(n10830), .B0(n8479), .B1(n7605), .Y(n10829)
         );
  OAI21X1 U9876 ( .A0(n12905), .A1(n7979), .B0(n8532), .Y(n10830) );
  AOI22X1 U9877 ( .A0(n8530), .A1(n8529), .B0(n12896), .B1(test_se), .Y(n10828) );
  NAND2X1 U9878 ( .A(n10831), .B(n10832), .Y(n6272) );
  AOI21X1 U9879 ( .A0(n10833), .A1(n8479), .B0(n10834), .Y(n10832) );
  AOI21X1 U9880 ( .A0(n8532), .A1(n10835), .B0(n7244), .Y(n10834) );
  NAND3X1 U9881 ( .A(n7944), .B(n7540), .C(n12490), .Y(n10835) );
  INVX1 U9882 ( .A(n8481), .Y(n8532) );
  NOR2X1 U9883 ( .A(n10836), .B(n7979), .Y(n8479) );
  INVX1 U9884 ( .A(n8480), .Y(n10833) );
  NAND3X1 U9885 ( .A(n10837), .B(n7244), .C(n12490), .Y(n8480) );
  AOI22X1 U9886 ( .A0(n7886), .A1(g29212), .B0(n12328), .B1(test_se), .Y(
        n10831) );
  OAI21X1 U9887 ( .A0(n7867), .A1(n7535), .B0(n10838), .Y(n6271) );
  AOI22X1 U9888 ( .A0(n12328), .A1(n10839), .B0(n12329), .B1(n8481), .Y(n10838) );
  OAI21X1 U9889 ( .A0(test_se), .A1(n10836), .B0(n7919), .Y(n10839) );
  INVX1 U9890 ( .A(n10840), .Y(n6270) );
  AOI22X1 U9891 ( .A0(n10841), .A1(n10842), .B0(n12329), .B1(n7979), .Y(n10840) );
  XOR2X1 U9892 ( .A(n12170), .B(n10843), .Y(n10842) );
  OAI21X1 U9893 ( .A0(n7944), .A1(n7696), .B0(n10844), .Y(n6269) );
  MX2X1 U9894 ( .A(n10845), .B(n10846), .S0(n7525), .Y(n10844) );
  NAND2X1 U9895 ( .A(n10847), .B(n10848), .Y(n10846) );
  NAND2X1 U9896 ( .A(n10841), .B(n10849), .Y(n10845) );
  OAI21X1 U9897 ( .A0(n7867), .A1(n7525), .B0(n10850), .Y(n6268) );
  AOI22X1 U9898 ( .A0(n12186), .A1(n8210), .B0(n12178), .B1(n8211), .Y(n10850)
         );
  NAND2X1 U9899 ( .A(n10851), .B(n10852), .Y(n6267) );
  AOI21X1 U9900 ( .A0(n8513), .A1(n7454), .B0(n10853), .Y(n10852) );
  AOI22X1 U9901 ( .A0(n12178), .A1(n7886), .B0(n12920), .B1(test_se), .Y(
        n10851) );
  NAND2X1 U9902 ( .A(n10854), .B(n10855), .Y(n6266) );
  MX2X1 U9903 ( .A(n7920), .B(n10856), .S0(n7219), .Y(n10855) );
  NAND4X1 U9904 ( .A(n12164), .B(n8514), .C(n12162), .D(n7357), .Y(n10856) );
  AOI21X1 U9905 ( .A0(test_se), .A1(n7454), .B0(n10857), .Y(n10854) );
  AOI21X1 U9906 ( .A0(n10858), .A1(n10859), .B0(n7407), .Y(n10857) );
  OAI21X1 U9907 ( .A0(n12165), .A1(n10860), .B0(n7923), .Y(n10859) );
  OAI21X1 U9908 ( .A0(n12160), .A1(n7867), .B0(n10861), .Y(n6265) );
  AOI21X1 U9909 ( .A0(n10862), .A1(n7296), .B0(n10863), .Y(n10861) );
  AOI21X1 U9910 ( .A0(n7921), .A1(n10864), .B0(n7407), .Y(n10863) );
  NAND3X1 U9911 ( .A(n10865), .B(n12166), .C(n12165), .Y(n10864) );
  NAND2X1 U9912 ( .A(n10858), .B(n10866), .Y(n10862) );
  NAND3X1 U9913 ( .A(n10867), .B(n10860), .C(n7944), .Y(n10866) );
  AOI21X1 U9914 ( .A0(n10868), .A1(n7944), .B0(n12165), .Y(n6264) );
  XOR2X1 U9915 ( .A(n7464), .B(n10869), .Y(n10868) );
  NOR2X1 U9916 ( .A(n10870), .B(n7219), .Y(n10869) );
  OAI21X1 U9917 ( .A0(n7867), .A1(n7464), .B0(n10871), .Y(n6263) );
  AOI22X1 U9918 ( .A0(n12489), .A1(n8559), .B0(n12166), .B1(n8513), .Y(n10871)
         );
  OAI21X1 U9919 ( .A0(n7867), .A1(n7573), .B0(n10872), .Y(n6262) );
  AOI21X1 U9920 ( .A0(n10873), .A1(n12167), .B0(n10874), .Y(n10872) );
  AOI21X1 U9921 ( .A0(n7920), .A1(n10875), .B0(n7464), .Y(n10874) );
  NAND4X1 U9922 ( .A(n10865), .B(n12166), .C(n7680), .D(n7296), .Y(n10875) );
  AOI21X1 U9923 ( .A0(n10858), .A1(n10876), .B0(n12165), .Y(n10873) );
  OAI21X1 U9924 ( .A0(n7219), .A1(n7464), .B0(n7922), .Y(n10876) );
  INVX1 U9925 ( .A(n8513), .Y(n10858) );
  OAI21X1 U9926 ( .A0(n8721), .A1(n7680), .B0(n10877), .Y(n6261) );
  AOI22X1 U9927 ( .A0(n10878), .A1(n12163), .B0(n10879), .B1(n8513), .Y(n10877) );
  NOR2X1 U9928 ( .A(n10880), .B(n10881), .Y(n10878) );
  NAND2X1 U9929 ( .A(n10882), .B(n10883), .Y(n6260) );
  MX2X1 U9930 ( .A(n10884), .B(n10885), .S0(n7368), .Y(n10883) );
  OR2X1 U9931 ( .A(n10886), .B(n10881), .Y(n10885) );
  AOI21X1 U9932 ( .A0(n12163), .A1(n7944), .B0(n8513), .Y(n10886) );
  NAND2X1 U9933 ( .A(n10879), .B(n10865), .Y(n10884) );
  AOI22X1 U9934 ( .A0(n7886), .A1(n7357), .B0(n12161), .B1(test_se), .Y(n10882) );
  NAND2X1 U9935 ( .A(n10887), .B(n10888), .Y(n6259) );
  MX2X1 U9936 ( .A(n10889), .B(n7867), .S0(n7357), .Y(n10888) );
  NAND3X1 U9937 ( .A(n12164), .B(n7944), .C(n10890), .Y(n10889) );
  AOI22X1 U9938 ( .A0(n10891), .A1(n10879), .B0(n7886), .B1(n7368), .Y(n10887)
         );
  NOR2X1 U9939 ( .A(n10892), .B(n9237), .Y(n10891) );
  XOR2X1 U9940 ( .A(n7461), .B(n10893), .Y(n10892) );
  NOR2X1 U9941 ( .A(n12160), .B(n10870), .Y(n10893) );
  OAI21X1 U9942 ( .A0(n8721), .A1(n7461), .B0(n10894), .Y(n6258) );
  MX2X1 U9943 ( .A(n10895), .B(n10896), .S0(n12161), .Y(n10894) );
  NAND2X1 U9944 ( .A(n10897), .B(n10890), .Y(n10896) );
  AOI21X1 U9945 ( .A0(n10898), .A1(n7357), .B0(n7979), .Y(n10897) );
  NAND2X1 U9946 ( .A(n10898), .B(n10879), .Y(n10895) );
  INVX1 U9947 ( .A(n10899), .Y(n10898) );
  NAND3X1 U9948 ( .A(n10900), .B(n7368), .C(n12164), .Y(n10899) );
  NAND2X1 U9949 ( .A(n10901), .B(n10902), .Y(n6257) );
  MX2X1 U9950 ( .A(n10903), .B(n10904), .S0(n7630), .Y(n10902) );
  NAND4X1 U9951 ( .A(n10905), .B(n10879), .C(n10865), .D(n12164), .Y(n10904)
         );
  NOR2X1 U9952 ( .A(n10881), .B(n12163), .Y(n10879) );
  NAND3X1 U9953 ( .A(n7944), .B(n10906), .C(n10890), .Y(n10903) );
  INVX1 U9954 ( .A(n10881), .Y(n10890) );
  OAI21X1 U9955 ( .A0(n7219), .A1(n7296), .B0(n10860), .Y(n10881) );
  NAND2X1 U9956 ( .A(n12167), .B(n12166), .Y(n10860) );
  NAND4X1 U9957 ( .A(n10905), .B(n12164), .C(n10900), .D(n7357), .Y(n10906) );
  INVX1 U9958 ( .A(n10867), .Y(n10905) );
  NAND2X1 U9959 ( .A(n12161), .B(n7368), .Y(n10867) );
  AOI22X1 U9960 ( .A0(n12161), .A1(n7885), .B0(test_se), .B1(n7251), .Y(n10901) );
  INVX1 U9961 ( .A(n10907), .Y(n6256) );
  AOI22X1 U9962 ( .A0(n10908), .A1(n7944), .B0(n12169), .B1(test_se), .Y(
        n10907) );
  XOR2X1 U9963 ( .A(n10909), .B(n10910), .Y(n10908) );
  XOR2X1 U9964 ( .A(n10911), .B(n10912), .Y(n10910) );
  XOR2X1 U9965 ( .A(n7206), .B(n10913), .Y(n10912) );
  NAND2X1 U9966 ( .A(n12159), .B(n10914), .Y(n10913) );
  XOR2X1 U9967 ( .A(n7397), .B(n7223), .Y(n10911) );
  XOR2X1 U9968 ( .A(n10915), .B(n10916), .Y(n10909) );
  XOR2X1 U9969 ( .A(n7222), .B(n7205), .Y(n10916) );
  XOR2X1 U9970 ( .A(n12938), .B(n7281), .Y(n10915) );
  NAND2X1 U9971 ( .A(n10917), .B(n10918), .Y(n6255) );
  MX2X1 U9972 ( .A(n12922), .B(n10919), .S0(n7870), .Y(n10918) );
  NAND2X1 U9973 ( .A(n10920), .B(n7619), .Y(n10919) );
  AOI22X1 U9974 ( .A0(n12225), .A1(n7885), .B0(n10921), .B1(n8562), .Y(n10917)
         );
  NOR2X1 U9975 ( .A(n10920), .B(n7619), .Y(n10921) );
  OAI21X1 U9976 ( .A0(n8721), .A1(n7619), .B0(n10922), .Y(n6254) );
  MX2X1 U9977 ( .A(n10923), .B(n12223), .S0(n10924), .Y(n10922) );
  NAND2X1 U9978 ( .A(n8562), .B(n12223), .Y(n10923) );
  OAI21X1 U9979 ( .A0(n7944), .A1(n7719), .B0(n10925), .Y(n6253) );
  MX2X1 U9980 ( .A(n10926), .B(n12222), .S0(n10927), .Y(n10925) );
  NAND2X1 U9981 ( .A(n8562), .B(n12222), .Y(n10926) );
  OAI21X1 U9982 ( .A0(n8721), .A1(n7720), .B0(n10928), .Y(n6252) );
  MX2X1 U9983 ( .A(n10929), .B(n12221), .S0(n10930), .Y(n10928) );
  NAND2X1 U9984 ( .A(n8562), .B(n12221), .Y(n10929) );
  OAI21X1 U9985 ( .A0(n7944), .A1(n7721), .B0(n10931), .Y(n6251) );
  MX2X1 U9986 ( .A(n10932), .B(n12220), .S0(n10933), .Y(n10931) );
  NAND2X1 U9987 ( .A(n8562), .B(n12220), .Y(n10932) );
  OAI21X1 U9988 ( .A0(n8721), .A1(n7722), .B0(n10934), .Y(n6250) );
  MX2X1 U9989 ( .A(n10935), .B(n12219), .S0(n10936), .Y(n10934) );
  NAND2X1 U9990 ( .A(n8562), .B(n12219), .Y(n10935) );
  OAI21X1 U9991 ( .A0(n7945), .A1(n7723), .B0(n10937), .Y(n6249) );
  MX2X1 U9992 ( .A(n10938), .B(n12218), .S0(n10939), .Y(n10937) );
  NAND2X1 U9993 ( .A(n8562), .B(n12218), .Y(n10938) );
  OAI21X1 U9994 ( .A0(n8721), .A1(n7724), .B0(n10940), .Y(n6248) );
  MX2X1 U9995 ( .A(n10941), .B(n12217), .S0(n10942), .Y(n10940) );
  NAND2X1 U9996 ( .A(n8562), .B(n12217), .Y(n10941) );
  OAI21X1 U9997 ( .A0(n7945), .A1(n7725), .B0(n10943), .Y(n6247) );
  MX2X1 U9998 ( .A(n10944), .B(n12228), .S0(n8644), .Y(n10943) );
  AND2X1 U9999 ( .A(n12217), .B(n10942), .Y(n8644) );
  AND2X1 U10000 ( .A(n12218), .B(n10939), .Y(n10942) );
  AND2X1 U10001 ( .A(n12219), .B(n10936), .Y(n10939) );
  AND2X1 U10002 ( .A(n12220), .B(n10933), .Y(n10936) );
  AND2X1 U10003 ( .A(n12221), .B(n10930), .Y(n10933) );
  AND2X1 U10004 ( .A(n12222), .B(n10927), .Y(n10930) );
  AND2X1 U10005 ( .A(n12223), .B(n10924), .Y(n10927) );
  AND2X1 U10006 ( .A(n12224), .B(n10920), .Y(n10924) );
  AND2X1 U10007 ( .A(n12225), .B(n10945), .Y(n10920) );
  NAND2X1 U10008 ( .A(n8562), .B(n12228), .Y(n10944) );
  OAI21X1 U10009 ( .A0(n7867), .A1(n7810), .B0(n10946), .Y(n6246) );
  AOI21X1 U10010 ( .A0(n12242), .A1(n7885), .B0(n10947), .Y(n10946) );
  AOI21X1 U10011 ( .A0(n12920), .A1(n7754), .B0(n10948), .Y(n10947) );
  OAI21X1 U10012 ( .A0(n7867), .A1(n7754), .B0(n10949), .Y(n6245) );
  AOI21X1 U10013 ( .A0(n12245), .A1(n7885), .B0(n10950), .Y(n10949) );
  AOI21X1 U10014 ( .A0(n12920), .A1(n7755), .B0(n7979), .Y(n10950) );
  OAI21X1 U10015 ( .A0(n7867), .A1(n7755), .B0(n10951), .Y(n6244) );
  AOI21X1 U10016 ( .A0(n12246), .A1(n7885), .B0(n10952), .Y(n10951) );
  AOI21X1 U10017 ( .A0(n7756), .A1(g29212), .B0(n7979), .Y(n10952) );
  OAI21X1 U10018 ( .A0(n7647), .A1(n7867), .B0(n10953), .Y(n6243) );
  AOI22X1 U10019 ( .A0(n12950), .A1(n7885), .B0(n7945), .B1(g21292), .Y(n10953) );
  NAND2X1 U10020 ( .A(n10954), .B(n10955), .Y(n6242) );
  MX2X1 U10021 ( .A(g30329), .B(n10956), .S0(n8104), .Y(n10955) );
  NAND2X1 U10022 ( .A(n8121), .B(n7681), .Y(n10956) );
  AOI22X1 U10023 ( .A0(n12915), .A1(n7885), .B0(n10957), .B1(n10958), .Y(
        n10954) );
  NOR2X1 U10024 ( .A(n8121), .B(n7681), .Y(n10957) );
  NOR2X1 U10025 ( .A(n7613), .B(n10959), .Y(n8121) );
  INVX1 U10026 ( .A(n10960), .Y(n6241) );
  AOI22X1 U10027 ( .A0(n8652), .A1(n10961), .B0(n12914), .B1(n7979), .Y(n10960) );
  XOR2X1 U10028 ( .A(n12904), .B(n10962), .Y(n10961) );
  NAND2X1 U10029 ( .A(n10963), .B(n10964), .Y(n6240) );
  MX2X1 U10030 ( .A(n12899), .B(n10965), .S0(n10966), .Y(n10964) );
  NAND2X1 U10031 ( .A(n12899), .B(n8652), .Y(n10965) );
  AOI22X1 U10032 ( .A0(n12900), .A1(n7885), .B0(n12904), .B1(test_se), .Y(
        n10963) );
  OAI21X1 U10033 ( .A0(n7945), .A1(n7682), .B0(n10967), .Y(n6239) );
  MX2X1 U10034 ( .A(n10968), .B(n12898), .S0(n10969), .Y(n10967) );
  NAND2X1 U10035 ( .A(n12898), .B(n8652), .Y(n10968) );
  OAI21X1 U10036 ( .A0(n8721), .A1(n7726), .B0(n10970), .Y(n6238) );
  MX2X1 U10037 ( .A(n10971), .B(n12894), .S0(n10972), .Y(n10970) );
  NAND2X1 U10038 ( .A(n12894), .B(n8652), .Y(n10971) );
  OAI21X1 U10039 ( .A0(n7945), .A1(n7727), .B0(n10973), .Y(n6237) );
  MX2X1 U10040 ( .A(n10974), .B(n10975), .S0(n7316), .Y(n10973) );
  NAND2X1 U10041 ( .A(n8652), .B(n10975), .Y(n10974) );
  NOR2X1 U10042 ( .A(n10976), .B(n7978), .Y(n8652) );
  OAI22X1 U10043 ( .A0(n7867), .A1(n7613), .B0(n10977), .B1(n7316), .Y(n6236)
         );
  AOI21X1 U10044 ( .A0(n10978), .A1(n7867), .B0(n7885), .Y(n10977) );
  INVX1 U10045 ( .A(n10975), .Y(n10978) );
  NAND2X1 U10046 ( .A(n12894), .B(n10972), .Y(n10975) );
  AND2X1 U10047 ( .A(n12898), .B(n10969), .Y(n10972) );
  NOR2X1 U10048 ( .A(n7682), .B(n10966), .Y(n10969) );
  NAND3X1 U10049 ( .A(n8649), .B(n8648), .C(n12900), .Y(n10966) );
  AND2X1 U10050 ( .A(n10962), .B(n12904), .Y(n8648) );
  INVX1 U10051 ( .A(n10976), .Y(n8649) );
  NAND3X1 U10052 ( .A(n10979), .B(n10980), .C(n12920), .Y(n10976) );
  OAI21X1 U10053 ( .A0(n12901), .A1(n10981), .B0(n10962), .Y(n10979) );
  INVX1 U10054 ( .A(n10982), .Y(n6235) );
  AOI22X1 U10055 ( .A0(g18099), .A1(n7945), .B0(n12777), .B1(test_se), .Y(
        n10982) );
  MX2X1 U10056 ( .A(g18098), .B(n13060), .S0(n7952), .Y(n6234) );
  OAI21X1 U10057 ( .A0(n7867), .A1(n7224), .B0(n10983), .Y(n6233) );
  AOI22X1 U10058 ( .A0(n10984), .A1(n7945), .B0(n13059), .B1(n7885), .Y(n10983) );
  MX2X1 U10059 ( .A(n10985), .B(n12590), .S0(n7956), .Y(n6232) );
  NAND2X1 U10060 ( .A(n7224), .B(n7207), .Y(n10985) );
  MX2X1 U10061 ( .A(n13059), .B(n7502), .S0(n8104), .Y(n6231) );
  INVX1 U10062 ( .A(n10986), .Y(n6230) );
  AOI21X1 U10063 ( .A0(n13057), .A1(n8593), .B0(n10987), .Y(n10986) );
  AOI21X1 U10064 ( .A0(n10988), .A1(n10989), .B0(n7978), .Y(n10987) );
  NAND4X1 U10065 ( .A(n12589), .B(n7207), .C(n7224), .D(n7811), .Y(n10989) );
  OAI21X1 U10066 ( .A0(n7502), .A1(n10990), .B0(n10984), .Y(n10988) );
  MX2X1 U10067 ( .A(n13060), .B(n13058), .S0(n7520), .Y(n10990) );
  OAI21X1 U10068 ( .A0(n7867), .A1(n7342), .B0(n10991), .Y(n6229) );
  AOI22X1 U10069 ( .A0(n7945), .A1(n10992), .B0(n13058), .B1(n7885), .Y(n10991) );
  OR2X1 U10070 ( .A(n10993), .B(n10994), .Y(n10992) );
  AOI21X1 U10071 ( .A0(n13058), .A1(n7283), .B0(n7520), .Y(n10994) );
  AOI21X1 U10072 ( .A0(n7224), .A1(n7283), .B0(n7207), .Y(n10993) );
  OAI21X1 U10073 ( .A0(n12589), .A1(n7867), .B0(n10995), .Y(n6228) );
  AOI22X1 U10074 ( .A0(n7945), .A1(n10996), .B0(n12588), .B1(n7885), .Y(n10995) );
  OAI21X1 U10075 ( .A0(n13058), .A1(n7283), .B0(n7207), .Y(n10996) );
  MX2X1 U10076 ( .A(n12532), .B(g8719), .S0(n8104), .Y(n6227) );
  MX2X1 U10077 ( .A(n10997), .B(n12931), .S0(n7953), .Y(n6226) );
  XOR2X1 U10078 ( .A(n12933), .B(n12934), .Y(n10997) );
  OAI21X1 U10079 ( .A0(n12932), .A1(n10998), .B0(n10999), .Y(n6225) );
  MX2X1 U10080 ( .A(n11000), .B(n7512), .S0(n7950), .Y(n10999) );
  NAND2X1 U10081 ( .A(n12932), .B(n10998), .Y(n11000) );
  OAI21X1 U10082 ( .A0(n5902), .A1(n7867), .B0(n11001), .Y(n6224) );
  AOI22X1 U10083 ( .A0(n7945), .A1(n11002), .B0(n7884), .B1(n12934), .Y(n11001) );
  XOR2X1 U10084 ( .A(n7536), .B(n8111), .Y(n11002) );
  NAND3X1 U10085 ( .A(n12932), .B(g8719), .C(n12933), .Y(n8111) );
  OAI21X1 U10086 ( .A0(n7867), .A1(n7812), .B0(n11003), .Y(n6223) );
  AOI22X1 U10087 ( .A0(n12439), .A1(n8559), .B0(n12476), .B1(n8513), .Y(n11003) );
  OAI21X1 U10088 ( .A0(n7867), .A1(n7728), .B0(n11004), .Y(n6222) );
  AOI22X1 U10089 ( .A0(n12435), .A1(n8559), .B0(n12439), .B1(n8513), .Y(n11004) );
  NAND2X1 U10090 ( .A(n11005), .B(n11006), .Y(n6221) );
  AOI22X1 U10091 ( .A0(n11007), .A1(n12850), .B0(n11008), .B1(n12772), .Y(
        n11006) );
  AOI22X1 U10092 ( .A0(n13066), .A1(n7884), .B0(n12439), .B1(test_se), .Y(
        n11005) );
  OAI21X1 U10093 ( .A0(n7867), .A1(n7575), .B0(n11009), .Y(n6220) );
  AOI22X1 U10094 ( .A0(n8513), .A1(n12477), .B0(n12850), .B1(n8514), .Y(n11009) );
  OAI21X1 U10095 ( .A0(n7866), .A1(n7370), .B0(n11010), .Y(n6219) );
  AOI22X1 U10096 ( .A0(n12478), .A1(n8559), .B0(n12475), .B1(n8513), .Y(n11010) );
  OAI21X1 U10097 ( .A0(n7866), .A1(n7373), .B0(n11011), .Y(n6218) );
  AOI22X1 U10098 ( .A0(n12487), .A1(n8559), .B0(n12491), .B1(n8513), .Y(n11011) );
  NAND2X1 U10099 ( .A(n11012), .B(n11013), .Y(n6217) );
  AOI22X1 U10100 ( .A0(n11014), .A1(n12489), .B0(n12488), .B1(n8513), .Y(
        n11013) );
  NOR2X1 U10101 ( .A(n12490), .B(n10880), .Y(n11014) );
  AOI22X1 U10102 ( .A0(n12491), .A1(n7884), .B0(n12932), .B1(test_se), .Y(
        n11012) );
  OAI21X1 U10103 ( .A0(n7866), .A1(n7729), .B0(n11015), .Y(n6216) );
  AOI22X1 U10104 ( .A0(n12488), .A1(n8559), .B0(n12851), .B1(n8513), .Y(n11015) );
  OR2X1 U10105 ( .A(n7884), .B(n10865), .Y(n8559) );
  NAND2X1 U10106 ( .A(n11016), .B(n11017), .Y(n6215) );
  AOI22X1 U10107 ( .A0(n11018), .A1(n12850), .B0(n12903), .B1(n8655), .Y(
        n11017) );
  NOR2X1 U10108 ( .A(n7978), .B(n11019), .Y(n11018) );
  AOI22X1 U10109 ( .A0(n12851), .A1(n7884), .B0(n12902), .B1(test_se), .Y(
        n11016) );
  MX2X1 U10110 ( .A(n12903), .B(g8358), .S0(n7847), .Y(n6214) );
  OAI21X1 U10111 ( .A0(n7866), .A1(n7631), .B0(n11020), .Y(n6213) );
  AOI22X1 U10112 ( .A0(n11021), .A1(n7945), .B0(n12827), .B1(n7884), .Y(n11020) );
  XOR2X1 U10113 ( .A(n11022), .B(n7800), .Y(n11021) );
  NAND2X1 U10114 ( .A(n11023), .B(n11024), .Y(n11022) );
  OAI21X1 U10115 ( .A0(n7866), .A1(n7841), .B0(n11025), .Y(n6212) );
  AOI22X1 U10116 ( .A0(n11026), .A1(n7945), .B0(n12828), .B1(n7884), .Y(n11025) );
  MX2X1 U10117 ( .A(n12892), .B(n11027), .S0(n11023), .Y(n11026) );
  NOR2X1 U10118 ( .A(n7828), .B(n12829), .Y(n11023) );
  INVX1 U10119 ( .A(n11024), .Y(n11027) );
  XOR2X1 U10120 ( .A(n7631), .B(g8358), .Y(n11024) );
  NAND2X1 U10121 ( .A(n11028), .B(n11029), .Y(n6211) );
  AOI22X1 U10122 ( .A0(n11007), .A1(n12940), .B0(n11008), .B1(g14189), .Y(
        n11029) );
  AOI22X1 U10123 ( .A0(n12772), .A1(n7884), .B0(n12827), .B1(test_se), .Y(
        n11028) );
  NAND2X1 U10124 ( .A(n11030), .B(n11031), .Y(n6210) );
  AOI22X1 U10125 ( .A0(n11007), .A1(n12935), .B0(n11008), .B1(g14201), .Y(
        n11031) );
  AOI22X1 U10126 ( .A0(n12940), .A1(n7884), .B0(n13066), .B1(test_se), .Y(
        n11030) );
  NAND2X1 U10127 ( .A(n11032), .B(n11033), .Y(n6209) );
  AOI22X1 U10128 ( .A0(n11007), .A1(n12937), .B0(n11008), .B1(g14217), .Y(
        n11033) );
  AOI22X1 U10129 ( .A0(n12935), .A1(n7884), .B0(n12940), .B1(test_se), .Y(
        n11032) );
  NAND2X1 U10130 ( .A(n11034), .B(n11035), .Y(n6208) );
  AOI22X1 U10131 ( .A0(n11007), .A1(n12938), .B0(n11008), .B1(g14096), .Y(
        n11035) );
  AOI22X1 U10132 ( .A0(n12937), .A1(n7884), .B0(n12935), .B1(test_se), .Y(
        n11034) );
  NAND2X1 U10133 ( .A(n11036), .B(n11037), .Y(n6207) );
  AOI22X1 U10134 ( .A0(n11007), .A1(n12939), .B0(n11008), .B1(g14125), .Y(
        n11037) );
  AOI22X1 U10135 ( .A0(n12938), .A1(n7884), .B0(n12937), .B1(test_se), .Y(
        n11036) );
  NAND2X1 U10136 ( .A(n11038), .B(n11039), .Y(n6206) );
  AOI22X1 U10137 ( .A0(n11007), .A1(n7205), .B0(n11008), .B1(g14147), .Y(
        n11039) );
  AOI22X1 U10138 ( .A0(n12939), .A1(n7883), .B0(n12938), .B1(test_se), .Y(
        n11038) );
  NAND2X1 U10139 ( .A(n11040), .B(n11041), .Y(n6205) );
  AOI22X1 U10140 ( .A0(n11007), .A1(n13066), .B0(n11008), .B1(g14167), .Y(
        n11041) );
  NOR2X1 U10141 ( .A(n11042), .B(n7978), .Y(n11008) );
  AND2X1 U10142 ( .A(n7945), .B(n11042), .Y(n11007) );
  NAND3X1 U10143 ( .A(n12771), .B(n7528), .C(n12770), .Y(n11042) );
  AOI22X1 U10144 ( .A0(n7883), .A1(n7205), .B0(n12939), .B1(test_se), .Y(
        n11040) );
  OAI21X1 U10145 ( .A0(n7538), .A1(n11043), .B0(n11044), .Y(n6204) );
  OAI21X1 U10146 ( .A0(n11045), .A1(test_se), .B0(n7205), .Y(n11044) );
  NOR2X1 U10147 ( .A(n11046), .B(n11047), .Y(n11045) );
  NAND3X1 U10148 ( .A(n12935), .B(n7945), .C(n12938), .Y(n11047) );
  NAND4X1 U10149 ( .A(n7206), .B(n7223), .C(n7397), .D(n7281), .Y(n11046) );
  OAI21X1 U10150 ( .A0(n11048), .A1(n11049), .B0(n7922), .Y(n11043) );
  NAND3X1 U10151 ( .A(n12937), .B(n12936), .C(n12940), .Y(n11049) );
  NAND4X1 U10152 ( .A(n12939), .B(n13066), .C(n7286), .D(n7222), .Y(n11048) );
  OAI22X1 U10153 ( .A0(n11050), .A1(n12919), .B0(n7538), .B1(n7945), .Y(n6203)
         );
  MX2X1 U10154 ( .A(n11051), .B(n11052), .S0(n12919), .Y(n6202) );
  OAI21X1 U10155 ( .A0(n11053), .A1(n7503), .B0(n8721), .Y(n11052) );
  NOR2X1 U10156 ( .A(n12918), .B(n11050), .Y(n11051) );
  OAI21X1 U10157 ( .A0(n12918), .A1(n7945), .B0(n11054), .Y(n6201) );
  MX2X1 U10158 ( .A(n12917), .B(n11055), .S0(n11056), .Y(n11054) );
  NAND2X1 U10159 ( .A(n10958), .B(n12917), .Y(n11055) );
  MX2X1 U10160 ( .A(n11057), .B(n11058), .S0(n12917), .Y(n6200) );
  NAND2X1 U10161 ( .A(n11059), .B(n8721), .Y(n11058) );
  MX2X1 U10162 ( .A(n12916), .B(n11060), .S0(n11056), .Y(n11059) );
  NAND2X1 U10163 ( .A(n12916), .B(n11061), .Y(n11060) );
  NOR2X1 U10164 ( .A(n7614), .B(n11050), .Y(n11057) );
  INVX1 U10165 ( .A(n10958), .Y(n11050) );
  OAI21X1 U10166 ( .A0(n7937), .A1(n7614), .B0(n11062), .Y(n6199) );
  MX2X1 U10167 ( .A(n12915), .B(n11063), .S0(n10959), .Y(n11062) );
  NAND3X1 U10168 ( .A(n12917), .B(n11064), .C(n12916), .Y(n10959) );
  INVX1 U10169 ( .A(n11056), .Y(n11064) );
  NAND3X1 U10170 ( .A(n11061), .B(n7503), .C(n12919), .Y(n11056) );
  INVX1 U10171 ( .A(n11053), .Y(n11061) );
  NAND2X1 U10172 ( .A(n10958), .B(n12915), .Y(n11063) );
  NOR2X1 U10173 ( .A(n11053), .B(n7978), .Y(n10958) );
  NAND4X1 U10174 ( .A(n12920), .B(n10980), .C(n11065), .D(n11066), .Y(n11053)
         );
  NOR2X1 U10175 ( .A(n11067), .B(n11068), .Y(n11066) );
  NAND2X1 U10176 ( .A(n11069), .B(n11070), .Y(n11068) );
  MX2X1 U10177 ( .A(n7222), .B(n7281), .S0(n7205), .Y(n11070) );
  MX2X1 U10178 ( .A(n12939), .B(n7538), .S0(n7223), .Y(n11069) );
  MX2X1 U10179 ( .A(n7222), .B(n7538), .S0(n7286), .Y(n11067) );
  MX2X1 U10180 ( .A(n12937), .B(n7397), .S0(n7206), .Y(n11065) );
  NAND2X1 U10181 ( .A(n11071), .B(n11072), .Y(n6198) );
  MX2X1 U10182 ( .A(n11073), .B(n11074), .S0(n7370), .Y(n11072) );
  OR2X1 U10183 ( .A(n10880), .B(n8668), .Y(n11074) );
  INVX1 U10184 ( .A(n8514), .Y(n10880) );
  AOI21X1 U10185 ( .A0(n10865), .A1(n8668), .B0(n7883), .Y(n11073) );
  XOR2X1 U10186 ( .A(n7370), .B(n11075), .Y(n8668) );
  AOI21X1 U10187 ( .A0(n12476), .A1(n11076), .B0(n11077), .Y(n11075) );
  MX2X1 U10188 ( .A(n11078), .B(n11079), .S0(n7373), .Y(n11077) );
  NOR2X1 U10189 ( .A(n12851), .B(n7321), .Y(n11079) );
  AND2X1 U10190 ( .A(n12851), .B(n12491), .Y(n11078) );
  XOR2X1 U10191 ( .A(n12488), .B(n12851), .Y(n11076) );
  NOR2X1 U10192 ( .A(n10870), .B(test_se), .Y(n10865) );
  AOI22X1 U10193 ( .A0(n12478), .A1(n8513), .B0(n12851), .B1(test_se), .Y(
        n11071) );
  OAI21X1 U10194 ( .A0(n7866), .A1(n7606), .B0(n11080), .Y(n6197) );
  AOI22X1 U10195 ( .A0(n12414), .A1(n8654), .B0(n12415), .B1(n8655), .Y(n11080) );
  OAI21X1 U10196 ( .A0(test_se), .A1(n11019), .B0(n7920), .Y(n8654) );
  NAND2X1 U10197 ( .A(n11081), .B(n11082), .Y(n6196) );
  AOI22X1 U10198 ( .A0(n11083), .A1(n11084), .B0(n12414), .B1(n8655), .Y(
        n11082) );
  NOR2X1 U10199 ( .A(n7978), .B(n11084), .Y(n8655) );
  NOR2X1 U10200 ( .A(n7978), .B(n7206), .Y(n11083) );
  AOI22X1 U10201 ( .A0(n12901), .A1(n7883), .B0(n12415), .B1(test_se), .Y(
        n11081) );
  NAND2X1 U10202 ( .A(n11085), .B(n11086), .Y(n6195) );
  AOI22X1 U10203 ( .A0(n12435), .A1(n8513), .B0(n8514), .B1(n13066), .Y(n11086) );
  NOR2X1 U10204 ( .A(n10870), .B(n7978), .Y(n8514) );
  NOR2X1 U10205 ( .A(n7978), .B(n10900), .Y(n8513) );
  INVX1 U10206 ( .A(n10870), .Y(n10900) );
  AOI22X1 U10207 ( .A0(n12475), .A1(n7883), .B0(n12414), .B1(test_se), .Y(
        n11085) );
  INVX1 U10208 ( .A(n11087), .Y(n6194) );
  AOI22X1 U10209 ( .A0(n12267), .A1(n11088), .B0(n12905), .B1(n8481), .Y(
        n11087) );
  INVX1 U10210 ( .A(n11089), .Y(n6193) );
  AOI22X1 U10211 ( .A0(n12905), .A1(n11088), .B0(n12927), .B1(n8481), .Y(
        n11089) );
  NOR2X1 U10212 ( .A(n7978), .B(n8529), .Y(n8481) );
  OAI21X1 U10213 ( .A0(n11090), .A1(n10836), .B0(n7922), .Y(n11088) );
  INVX1 U10214 ( .A(n11091), .Y(n6192) );
  AOI22X1 U10215 ( .A0(n11092), .A1(n10962), .B0(n12435), .B1(test_se), .Y(
        n11091) );
  INVX1 U10216 ( .A(n11093), .Y(n10962) );
  NAND3X1 U10217 ( .A(n12927), .B(n7615), .C(n12906), .Y(n11093) );
  NOR2X1 U10218 ( .A(n11094), .B(n7978), .Y(n11092) );
  AOI22X1 U10219 ( .A0(n12901), .A1(n10981), .B0(n12903), .B1(n12902), .Y(
        n11094) );
  OR2X1 U10220 ( .A(n12902), .B(n12903), .Y(n10981) );
  AND2X1 U10221 ( .A(n11095), .B(n11096), .Y(n6191) );
  MX2X1 U10222 ( .A(n11097), .B(n12927), .S0(n7950), .Y(n11095) );
  MX2X1 U10223 ( .A(n11098), .B(n11099), .S0(n7284), .Y(n11097) );
  AOI21X1 U10224 ( .A0(n12929), .A1(n7365), .B0(n11098), .Y(n11099) );
  NAND2X1 U10225 ( .A(n11100), .B(n11101), .Y(n6190) );
  AOI21X1 U10226 ( .A0(n11102), .A1(n7934), .B0(n8530), .Y(n11101) );
  XOR2X1 U10227 ( .A(n7365), .B(n11103), .Y(n11102) );
  AOI22X1 U10228 ( .A0(n12930), .A1(n7883), .B0(test_se), .B1(n7460), .Y(
        n11100) );
  NAND2X1 U10229 ( .A(n11104), .B(n11105), .Y(n6189) );
  MX2X1 U10230 ( .A(n11106), .B(n12928), .S0(n7949), .Y(n11105) );
  NAND2X1 U10231 ( .A(n12929), .B(n11107), .Y(n11106) );
  AOI21X1 U10232 ( .A0(n11108), .A1(n7462), .B0(n8530), .Y(n11104) );
  INVX1 U10233 ( .A(n11096), .Y(n8530) );
  NAND2X1 U10234 ( .A(n11090), .B(n7934), .Y(n11096) );
  NOR2X1 U10235 ( .A(n7814), .B(n12328), .Y(n11090) );
  INVX1 U10236 ( .A(n11107), .Y(n11108) );
  NAND2X1 U10237 ( .A(n11103), .B(n7365), .Y(n11107) );
  NOR2X1 U10238 ( .A(n11109), .B(n11098), .Y(n11103) );
  NAND3X1 U10239 ( .A(n8529), .B(n7615), .C(n12927), .Y(n11098) );
  INVX1 U10240 ( .A(n10836), .Y(n8529) );
  NAND3X1 U10241 ( .A(n12934), .B(n7512), .C(n12932), .Y(n10836) );
  AOI21X1 U10242 ( .A0(n12929), .A1(n7365), .B0(n12930), .Y(n11109) );
  OAI21X1 U10243 ( .A0(n7866), .A1(n7284), .B0(n11110), .Y(n6188) );
  AOI21X1 U10244 ( .A0(n12247), .A1(n7883), .B0(n11111), .Y(n11110) );
  AOI21X1 U10245 ( .A0(n7757), .A1(n7343), .B0(n7978), .Y(n11111) );
  NAND2X1 U10246 ( .A(n11112), .B(n11113), .Y(n6187) );
  MX2X1 U10247 ( .A(n11114), .B(n11115), .S0(n12158), .Y(n11113) );
  AOI22X1 U10248 ( .A0(n12585), .A1(n7935), .B0(n12532), .B1(n7866), .Y(n11115) );
  NAND2X1 U10249 ( .A(n7935), .B(g29211), .Y(n11114) );
  AOI22X1 U10250 ( .A0(n12532), .A1(n7883), .B0(test_se), .B1(g18881), .Y(
        n11112) );
  NAND3X1 U10251 ( .A(n11116), .B(n11117), .C(n11118), .Y(n6186) );
  NAND2X1 U10252 ( .A(test_se), .B(g29215), .Y(n11118) );
  NAND4X1 U10253 ( .A(n13057), .B(n7935), .C(n11119), .D(n7820), .Y(n11117) );
  INVX1 U10254 ( .A(n10984), .Y(n11119) );
  MX2X1 U10255 ( .A(n13060), .B(n13058), .S0(n7283), .Y(n10984) );
  NAND2X1 U10256 ( .A(n7883), .B(g29211), .Y(n11116) );
  OAI21X1 U10257 ( .A0(n7866), .A1(n7520), .B0(n11120), .Y(n6185) );
  AOI22X1 U10258 ( .A0(n7883), .A1(g21176), .B0(n12590), .B1(n7935), .Y(n11120) );
  OAI21X1 U10259 ( .A0(n7866), .A1(n7820), .B0(n11121), .Y(n6184) );
  AOI22X1 U10260 ( .A0(n12585), .A1(n7883), .B0(n7935), .B1(n7661), .Y(n11121)
         );
  MX2X1 U10261 ( .A(n7977), .B(n11122), .S0(n7661), .Y(n6183) );
  NOR2X1 U10262 ( .A(n12533), .B(n7977), .Y(n11122) );
  NAND2X1 U10263 ( .A(n11123), .B(n11124), .Y(n6182) );
  AOI22X1 U10264 ( .A0(n9960), .A1(n9968), .B0(n10100), .B1(g21245), .Y(n11124) );
  NOR2X1 U10265 ( .A(n7977), .B(g33959), .Y(n10100) );
  NOR2X1 U10266 ( .A(n9987), .B(n7977), .Y(n9968) );
  MX2X1 U10267 ( .A(n11125), .B(n11126), .S0(g25219), .Y(n9960) );
  NAND4X1 U10268 ( .A(n11127), .B(n11128), .C(n11129), .D(n11130), .Y(n11126)
         );
  OR2X1 U10269 ( .A(n11131), .B(n10113), .Y(n11130) );
  AOI22X1 U10270 ( .A0(n12975), .A1(g13039), .B0(n12976), .B1(n12980), .Y(
        n11131) );
  AOI22X1 U10271 ( .A0(n11132), .A1(n12978), .B0(n11133), .B1(n12977), .Y(
        n11129) );
  NOR2X1 U10272 ( .A(n5261), .B(n10104), .Y(n11133) );
  NOR2X1 U10273 ( .A(n5260), .B(n10112), .Y(n11132) );
  OR2X1 U10274 ( .A(n11134), .B(n10114), .Y(n11128) );
  AOI22X1 U10275 ( .A0(g17639), .A1(n7227), .B0(n13005), .B1(g17577), .Y(
        n11134) );
  MX2X1 U10276 ( .A(n11135), .B(n11136), .S0(g12238), .Y(n11127) );
  AOI21X1 U10277 ( .A0(n11137), .A1(n7446), .B0(n11138), .Y(n11136) );
  INVX1 U10278 ( .A(n11139), .Y(n11135) );
  NAND4X1 U10279 ( .A(n11140), .B(n11141), .C(n11142), .D(n11143), .Y(n11125)
         );
  OR2X1 U10280 ( .A(n11144), .B(n10112), .Y(n11143) );
  AOI22X1 U10281 ( .A0(n12979), .A1(g13039), .B0(n12980), .B1(n12981), .Y(
        n11144) );
  AOI22X1 U10282 ( .A0(n11145), .A1(n12991), .B0(n11146), .B1(n12994), .Y(
        n11142) );
  NOR2X1 U10283 ( .A(n5261), .B(n10114), .Y(n11146) );
  NOR2X1 U10284 ( .A(n5260), .B(n10113), .Y(n11145) );
  INVX1 U10285 ( .A(n11147), .Y(n10113) );
  OR2X1 U10286 ( .A(n11148), .B(n10104), .Y(n11141) );
  INVX1 U10287 ( .A(n11137), .Y(n10104) );
  AOI22X1 U10288 ( .A0(n12990), .A1(g17639), .B0(n12989), .B1(g17577), .Y(
        n11148) );
  MX2X1 U10289 ( .A(n11149), .B(n11150), .S0(g12238), .Y(n11140) );
  AOI21X1 U10290 ( .A0(n12985), .A1(g25114), .B0(n11139), .Y(n11150) );
  NAND3X1 U10291 ( .A(n11151), .B(n11152), .C(n11153), .Y(n11139) );
  NAND3X1 U10292 ( .A(n11147), .B(g14662), .C(n12982), .Y(n11153) );
  NAND3X1 U10293 ( .A(n10101), .B(g17519), .C(n12984), .Y(n11152) );
  NAND3X1 U10294 ( .A(n11137), .B(g17674), .C(n12983), .Y(n11151) );
  NOR2X1 U10295 ( .A(n12993), .B(n12992), .Y(n11137) );
  INVX1 U10296 ( .A(n11138), .Y(n11149) );
  NAND3X1 U10297 ( .A(n11154), .B(n11155), .C(n11156), .Y(n11138) );
  NAND3X1 U10298 ( .A(g25114), .B(g17674), .C(n12986), .Y(n11156) );
  NAND3X1 U10299 ( .A(n10101), .B(g14662), .C(n12987), .Y(n11155) );
  INVX1 U10300 ( .A(n10112), .Y(n10101) );
  NAND2X1 U10301 ( .A(n12992), .B(n12993), .Y(n10112) );
  NAND3X1 U10302 ( .A(n11147), .B(g17519), .C(n12988), .Y(n11154) );
  NOR2X1 U10303 ( .A(n7366), .B(n12993), .Y(n11147) );
  AOI22X1 U10304 ( .A0(n13005), .A1(n7883), .B0(test_se), .B1(g29219), .Y(
        n11123) );
  NAND2X1 U10305 ( .A(n11157), .B(n11158), .Y(n6181) );
  AOI22X1 U10306 ( .A0(n11159), .A1(n7730), .B0(n11160), .B1(n7302), .Y(n11158) );
  AOI22X1 U10307 ( .A0(n7882), .A1(g29219), .B0(n12698), .B1(test_se), .Y(
        n11157) );
  OAI21X1 U10308 ( .A0(n12697), .A1(n7866), .B0(n11161), .Y(n6180) );
  AOI22X1 U10309 ( .A0(n11162), .A1(n7935), .B0(n7882), .B1(n7378), .Y(n11161)
         );
  MX2X1 U10310 ( .A(n7381), .B(n12697), .S0(n11163), .Y(n11162) );
  OAI21X1 U10311 ( .A0(n13020), .A1(n7866), .B0(n11164), .Y(n6179) );
  AOI22X1 U10312 ( .A0(n11165), .A1(n7935), .B0(n7882), .B1(n7271), .Y(n11164)
         );
  MX2X1 U10313 ( .A(n12688), .B(n7378), .S0(n11166), .Y(n11165) );
  NAND2X1 U10314 ( .A(n11167), .B(n11168), .Y(n6178) );
  AOI22X1 U10315 ( .A0(n11159), .A1(n7731), .B0(n11160), .B1(n7305), .Y(n11168) );
  AOI22X1 U10316 ( .A0(n7882), .A1(n7302), .B0(test_se), .B1(n7378), .Y(n11167) );
  OAI21X1 U10317 ( .A0(n12688), .A1(n7866), .B0(n11169), .Y(n6177) );
  AOI22X1 U10318 ( .A0(n11170), .A1(n7935), .B0(n7882), .B1(n7218), .Y(n11169)
         );
  MX2X1 U10319 ( .A(n7271), .B(n12687), .S0(n11171), .Y(n11170) );
  OAI21X1 U10320 ( .A0(n13021), .A1(n7866), .B0(n11172), .Y(n6176) );
  AOI22X1 U10321 ( .A0(n11173), .A1(n7935), .B0(n7882), .B1(n7306), .Y(n11172)
         );
  MX2X1 U10322 ( .A(n7218), .B(n12686), .S0(n11174), .Y(n11173) );
  NAND2X1 U10323 ( .A(n11175), .B(n11176), .Y(n6175) );
  AOI22X1 U10324 ( .A0(n11177), .A1(n11178), .B0(n12711), .B1(n11179), .Y(
        n11176) );
  NOR2X1 U10325 ( .A(n12710), .B(n11180), .Y(n11177) );
  AOI22X1 U10326 ( .A0(n12713), .A1(n7882), .B0(test_se), .B1(n7450), .Y(
        n11175) );
  NAND3X1 U10327 ( .A(n11181), .B(n11182), .C(n11183), .Y(n6174) );
  AOI22X1 U10328 ( .A0(n12710), .A1(n7882), .B0(n12722), .B1(test_se), .Y(
        n11183) );
  NAND2X1 U10329 ( .A(n11179), .B(n13023), .Y(n11182) );
  AOI22X1 U10330 ( .A0(n11184), .A1(n11185), .B0(n11178), .B1(n11186), .Y(
        n11181) );
  NAND3X1 U10331 ( .A(n11187), .B(n11188), .C(n11189), .Y(n11186) );
  AOI22X1 U10332 ( .A0(n11180), .A1(n7393), .B0(n12719), .B1(n11190), .Y(
        n11189) );
  NAND3X1 U10333 ( .A(n7487), .B(n7289), .C(n12715), .Y(n11188) );
  OR2X1 U10334 ( .A(n12712), .B(n11191), .Y(n11187) );
  AOI22X1 U10335 ( .A0(n12710), .A1(n12717), .B0(n12716), .B1(n12711), .Y(
        n11191) );
  INVX1 U10336 ( .A(n11192), .Y(n11185) );
  NOR2X1 U10337 ( .A(n12714), .B(n7977), .Y(n11184) );
  NAND2X1 U10338 ( .A(n11193), .B(n11194), .Y(n6173) );
  MX2X1 U10339 ( .A(n11195), .B(n11196), .S0(n7325), .Y(n11194) );
  NAND2X1 U10340 ( .A(n11197), .B(n7935), .Y(n11196) );
  AOI21X1 U10341 ( .A0(n11198), .A1(n8717), .B0(n7882), .Y(n11195) );
  NOR2X1 U10342 ( .A(n11199), .B(n11197), .Y(n11198) );
  NOR2X1 U10343 ( .A(n12706), .B(n11180), .Y(n11197) );
  AOI22X1 U10344 ( .A0(n11179), .A1(n7435), .B0(n12718), .B1(test_se), .Y(
        n11193) );
  OAI21X1 U10345 ( .A0(n12706), .A1(n8721), .B0(n11200), .Y(n6172) );
  AOI22X1 U10346 ( .A0(n11201), .A1(n11202), .B0(n12705), .B1(n11203), .Y(
        n11200) );
  OAI21X1 U10347 ( .A0(n11180), .A1(n7977), .B0(n11204), .Y(n11203) );
  INVX1 U10348 ( .A(n11179), .Y(n11204) );
  XOR2X1 U10349 ( .A(n12718), .B(n7435), .Y(n11202) );
  AND2X1 U10350 ( .A(n11178), .B(n11180), .Y(n11201) );
  NOR2X1 U10351 ( .A(n7553), .B(n12711), .Y(n11180) );
  OAI21X1 U10352 ( .A0(n7935), .A1(n7216), .B0(n11205), .Y(n6171) );
  MX2X1 U10353 ( .A(n11206), .B(n11207), .S0(n7586), .Y(n11205) );
  NAND2X1 U10354 ( .A(n11190), .B(n11178), .Y(n11207) );
  MX2X1 U10355 ( .A(n12703), .B(n12704), .S0(n11208), .Y(n6170) );
  OAI21X1 U10356 ( .A0(n11208), .A1(n7238), .B0(n11209), .Y(n6169) );
  MX2X1 U10357 ( .A(n11210), .B(n11211), .S0(n12703), .Y(n11209) );
  AOI21X1 U10358 ( .A0(n8373), .A1(n12704), .B0(n8593), .Y(n11211) );
  NAND3X1 U10359 ( .A(n7935), .B(n7586), .C(n8373), .Y(n11210) );
  OAI21X1 U10360 ( .A0(n11208), .A1(n7308), .B0(n11212), .Y(n6168) );
  MX2X1 U10361 ( .A(n11213), .B(n7238), .S0(n7952), .Y(n11212) );
  NAND2X1 U10362 ( .A(n8373), .B(n7308), .Y(n11213) );
  OAI22X1 U10363 ( .A0(n11206), .A1(n7662), .B0(n11214), .B1(n7308), .Y(n6167)
         );
  AOI21X1 U10364 ( .A0(n11190), .A1(n11215), .B0(n8593), .Y(n11214) );
  OAI21X1 U10365 ( .A0(n11206), .A1(n7213), .B0(n11216), .Y(n6166) );
  MX2X1 U10366 ( .A(n11217), .B(n11218), .S0(n7662), .Y(n11216) );
  NAND3X1 U10367 ( .A(n11178), .B(n7308), .C(n11190), .Y(n11218) );
  AOI21X1 U10368 ( .A0(n11219), .A1(n12702), .B0(n8593), .Y(n11217) );
  NOR2X1 U10369 ( .A(n11220), .B(n11221), .Y(n11219) );
  AOI21X1 U10370 ( .A0(n11221), .A1(n7935), .B0(n11179), .Y(n11206) );
  INVX1 U10371 ( .A(n11190), .Y(n11221) );
  NOR2X1 U10372 ( .A(n7289), .B(n7487), .Y(n11190) );
  OAI21X1 U10373 ( .A0(n7866), .A1(n7213), .B0(n7951), .Y(n6165) );
  NAND2X1 U10374 ( .A(n7320), .B(n7977), .Y(n6164) );
  NOR2X1 U10375 ( .A(n8721), .B(n7574), .Y(n6163) );
  NAND2X1 U10376 ( .A(n7492), .B(n7977), .Y(n6162) );
  NAND2X1 U10377 ( .A(n7300), .B(n7977), .Y(n6161) );
  NOR2X1 U10378 ( .A(n8721), .B(n7688), .Y(n6160) );
  NOR2X1 U10379 ( .A(n8721), .B(n7319), .Y(n6159) );
  OR2X1 U10380 ( .A(n13029), .B(n7935), .Y(n6158) );
  OAI21X1 U10381 ( .A0(n7866), .A1(n7457), .B0(n11222), .Y(n6157) );
  AOI22X1 U10382 ( .A0(n11223), .A1(n7935), .B0(n12785), .B1(n7882), .Y(n11222) );
  MX2X1 U10383 ( .A(n11224), .B(n12783), .S0(n11225), .Y(n11223) );
  NAND2X1 U10384 ( .A(n12791), .B(n7265), .Y(n11224) );
  NAND2X1 U10385 ( .A(n11226), .B(n11227), .Y(n6156) );
  AOI22X1 U10386 ( .A0(n11228), .A1(n12792), .B0(n8405), .B1(n12791), .Y(
        n11227) );
  NOR2X1 U10387 ( .A(n8413), .B(n7977), .Y(n11228) );
  AOI22X1 U10388 ( .A0(n12779), .A1(n7882), .B0(n12783), .B1(test_se), .Y(
        n11226) );
  OAI21X1 U10389 ( .A0(n7866), .A1(n7693), .B0(n11229), .Y(n6155) );
  AOI22X1 U10390 ( .A0(n12782), .A1(n11230), .B0(n8760), .B1(n12781), .Y(
        n11229) );
  OAI21X1 U10391 ( .A0(test_se), .A1(n11231), .B0(n7919), .Y(n11230) );
  OAI21X1 U10392 ( .A0(n7920), .A1(n7234), .B0(n11232), .Y(n6154) );
  AOI21X1 U10393 ( .A0(n8760), .A1(n12780), .B0(n11233), .Y(n11232) );
  AOI21X1 U10394 ( .A0(n7866), .A1(n11234), .B0(n7488), .Y(n11233) );
  INVX1 U10395 ( .A(n8766), .Y(n11234) );
  NAND2X1 U10396 ( .A(n11235), .B(n11236), .Y(n6153) );
  MX2X1 U10397 ( .A(n7234), .B(n11237), .S0(n7853), .Y(n11236) );
  AOI22X1 U10398 ( .A0(n12793), .A1(n8405), .B0(n12791), .B1(n7882), .Y(n11235) );
  NOR2X1 U10399 ( .A(n8749), .B(n7977), .Y(n8405) );
  NAND2X1 U10400 ( .A(n11238), .B(n11239), .Y(n6152) );
  AOI22X1 U10401 ( .A0(n11240), .A1(n11241), .B0(n12789), .B1(n11242), .Y(
        n11239) );
  AOI22X1 U10402 ( .A0(n12788), .A1(n7880), .B0(n12790), .B1(test_se), .Y(
        n11238) );
  NAND2X1 U10403 ( .A(n11243), .B(n11244), .Y(n6151) );
  MX2X1 U10404 ( .A(n11245), .B(n11246), .S0(n11247), .Y(n11244) );
  NOR2X1 U10405 ( .A(n7265), .B(n11248), .Y(n11247) );
  NAND2X1 U10406 ( .A(n8749), .B(n7465), .Y(n11248) );
  OAI21X1 U10407 ( .A0(n12893), .A1(n8414), .B0(g35), .Y(n11246) );
  NAND2X1 U10408 ( .A(n12790), .B(n7935), .Y(n11245) );
  AOI22X1 U10409 ( .A0(n12789), .A1(n7880), .B0(n12792), .B1(test_se), .Y(
        n11243) );
  NAND2X1 U10410 ( .A(n11249), .B(n11250), .Y(n6150) );
  MX2X1 U10411 ( .A(n11251), .B(n11252), .S0(n11253), .Y(n11250) );
  NOR2X1 U10412 ( .A(n12793), .B(n11237), .Y(n11253) );
  NAND2X1 U10413 ( .A(n12787), .B(n7935), .Y(n11251) );
  AOI22X1 U10414 ( .A0(n12790), .A1(n7880), .B0(n12789), .B1(test_se), .Y(
        n11249) );
  NAND2X1 U10415 ( .A(n11254), .B(n11255), .Y(n6149) );
  MX2X1 U10416 ( .A(n11256), .B(n11252), .S0(n11257), .Y(n11255) );
  NOR2X1 U10417 ( .A(n7265), .B(n8750), .Y(n11257) );
  NAND2X1 U10418 ( .A(n12785), .B(n7935), .Y(n11256) );
  AOI22X1 U10419 ( .A0(n12786), .A1(n7880), .B0(n12787), .B1(test_se), .Y(
        n11254) );
  NAND2X1 U10420 ( .A(n11258), .B(n11259), .Y(n6148) );
  MX2X1 U10421 ( .A(n11260), .B(n11252), .S0(n11261), .Y(n11259) );
  NOR2X1 U10422 ( .A(n12792), .B(n11237), .Y(n11261) );
  NAND2X1 U10423 ( .A(n12791), .B(n8749), .Y(n11237) );
  NAND2X1 U10424 ( .A(n12786), .B(n7935), .Y(n11260) );
  AOI22X1 U10425 ( .A0(n7880), .A1(n7447), .B0(n12785), .B1(test_se), .Y(
        n11258) );
  NAND2X1 U10426 ( .A(n11262), .B(n11263), .Y(n6147) );
  MX2X1 U10427 ( .A(n11264), .B(n11252), .S0(n11265), .Y(n11263) );
  NOR2X1 U10428 ( .A(n12791), .B(n8750), .Y(n11265) );
  NAND2X1 U10429 ( .A(n12793), .B(n8749), .Y(n8750) );
  INVX1 U10430 ( .A(n11240), .Y(n11252) );
  AOI21X1 U10431 ( .A0(n7474), .A1(n11266), .B0(n7977), .Y(n11240) );
  NAND2X1 U10432 ( .A(n7935), .B(n7447), .Y(n11264) );
  AOI22X1 U10433 ( .A0(n12787), .A1(n7880), .B0(n12786), .B1(test_se), .Y(
        n11262) );
  NAND2X1 U10434 ( .A(n11267), .B(n11268), .Y(n6146) );
  AOI21X1 U10435 ( .A0(n12782), .A1(n8760), .B0(n11269), .Y(n11268) );
  NOR2X1 U10436 ( .A(n12780), .B(n11270), .Y(n11269) );
  AOI22X1 U10437 ( .A0(n8766), .A1(n7488), .B0(n12782), .B1(n7935), .Y(n11270)
         );
  AOI22X1 U10438 ( .A0(n12783), .A1(n7880), .B0(test_se), .B1(n7447), .Y(
        n11267) );
  OAI21X1 U10439 ( .A0(n7935), .A1(n7765), .B0(n11271), .Y(n6145) );
  MX2X1 U10440 ( .A(n11272), .B(n11273), .S0(n7587), .Y(n11271) );
  NAND2X1 U10441 ( .A(n11274), .B(n8766), .Y(n11273) );
  MX2X1 U10442 ( .A(n12768), .B(n12773), .S0(n8751), .Y(n6144) );
  OAI21X1 U10443 ( .A0(n8751), .A1(n7763), .B0(n11275), .Y(n6143) );
  MX2X1 U10444 ( .A(n11276), .B(n11277), .S0(n12768), .Y(n11275) );
  AOI21X1 U10445 ( .A0(n12773), .A1(n11241), .B0(n8593), .Y(n11277) );
  NAND2X1 U10446 ( .A(n8411), .B(n7587), .Y(n11276) );
  INVX1 U10447 ( .A(n11242), .Y(n8751) );
  INVX1 U10448 ( .A(n11278), .Y(n6142) );
  AOI21X1 U10449 ( .A0(n7977), .A1(n12767), .B0(n11279), .Y(n11278) );
  MX2X1 U10450 ( .A(n11242), .B(n8411), .S0(n7521), .Y(n11279) );
  NOR2X1 U10451 ( .A(n11280), .B(n7976), .Y(n8411) );
  NOR2X1 U10452 ( .A(n7976), .B(n11241), .Y(n11242) );
  INVX1 U10453 ( .A(n11280), .Y(n11241) );
  NAND3X1 U10454 ( .A(n7497), .B(n7265), .C(n8749), .Y(n11280) );
  INVX1 U10455 ( .A(n8413), .Y(n8749) );
  NOR2X1 U10456 ( .A(n11281), .B(n8414), .Y(n8413) );
  INVX1 U10457 ( .A(n11266), .Y(n8414) );
  NOR2X1 U10458 ( .A(n11282), .B(n12913), .Y(n11266) );
  AOI21X1 U10459 ( .A0(n10694), .A1(n11283), .B0(n5266), .Y(n11281) );
  INVX1 U10460 ( .A(n10782), .Y(n10694) );
  NAND2X1 U10461 ( .A(n12973), .B(n7551), .Y(n10782) );
  OAI21X1 U10462 ( .A0(n8721), .A1(n7521), .B0(n11284), .Y(n6141) );
  AOI21X1 U10463 ( .A0(n12765), .A1(n11285), .B0(n11286), .Y(n11284) );
  OAI21X1 U10464 ( .A0(n11272), .A1(n7335), .B0(n11287), .Y(n6140) );
  MX2X1 U10465 ( .A(n11288), .B(n11289), .S0(n12765), .Y(n11287) );
  NOR2X1 U10466 ( .A(n11286), .B(n8593), .Y(n11289) );
  INVX1 U10467 ( .A(n11290), .Y(n11286) );
  NAND3X1 U10468 ( .A(n11274), .B(n8758), .C(n12766), .Y(n11290) );
  NAND3X1 U10469 ( .A(n8766), .B(n7521), .C(n11274), .Y(n11288) );
  INVX1 U10470 ( .A(n11285), .Y(n11272) );
  OAI21X1 U10471 ( .A0(n11274), .A1(n7976), .B0(n8765), .Y(n11285) );
  INVX1 U10472 ( .A(n8760), .Y(n8765) );
  OAI22X1 U10473 ( .A0(n7866), .A1(n7335), .B0(n11291), .B1(n7976), .Y(n6139)
         );
  AOI22X1 U10474 ( .A0(n11292), .A1(n11293), .B0(n12763), .B1(n11294), .Y(
        n11291) );
  NOR2X1 U10475 ( .A(n12762), .B(n12764), .Y(n11292) );
  MX2X1 U10476 ( .A(n12760), .B(n12749), .S0(n11295), .Y(n6138) );
  NAND2X1 U10477 ( .A(n11296), .B(n11297), .Y(n6137) );
  AOI22X1 U10478 ( .A0(n11298), .A1(n8399), .B0(n12761), .B1(n11299), .Y(
        n11297) );
  INVX1 U10479 ( .A(n11300), .Y(n11298) );
  AOI22X1 U10480 ( .A0(n12760), .A1(n7880), .B0(test_se), .B1(n7391), .Y(
        n11296) );
  NAND2X1 U10481 ( .A(n11301), .B(n11302), .Y(n6136) );
  MX2X1 U10482 ( .A(n11303), .B(n11300), .S0(n11304), .Y(n11302) );
  NOR2X1 U10483 ( .A(n12764), .B(n11305), .Y(n11304) );
  NAND2X1 U10484 ( .A(n12759), .B(n7935), .Y(n11303) );
  AOI22X1 U10485 ( .A0(n7880), .A1(n7391), .B0(n12761), .B1(test_se), .Y(
        n11301) );
  NAND2X1 U10486 ( .A(n11306), .B(n11307), .Y(n6135) );
  MX2X1 U10487 ( .A(n11308), .B(n11300), .S0(n11309), .Y(n11307) );
  NOR2X1 U10488 ( .A(n12762), .B(n11294), .Y(n11309) );
  NAND2X1 U10489 ( .A(n7935), .B(n7448), .Y(n11308) );
  AOI22X1 U10490 ( .A0(n12759), .A1(n7880), .B0(n12758), .B1(test_se), .Y(
        n11306) );
  NAND2X1 U10491 ( .A(n11310), .B(n11311), .Y(n6134) );
  AOI22X1 U10492 ( .A0(n11312), .A1(n11313), .B0(n12753), .B1(n11314), .Y(
        n11311) );
  NOR2X1 U10493 ( .A(n12752), .B(n11315), .Y(n11312) );
  AOI22X1 U10494 ( .A0(n12755), .A1(n7880), .B0(test_se), .B1(n7448), .Y(
        n11310) );
  OAI21X1 U10495 ( .A0(n7866), .A1(n7485), .B0(n11316), .Y(n6133) );
  AOI22X1 U10496 ( .A0(n11317), .A1(n7936), .B0(n12757), .B1(n7880), .Y(n11316) );
  MX2X1 U10497 ( .A(n11318), .B(n12755), .S0(n11319), .Y(n11317) );
  NAND2X1 U10498 ( .A(n12762), .B(n7400), .Y(n11318) );
  NAND2X1 U10499 ( .A(n11320), .B(n11321), .Y(n6132) );
  AOI22X1 U10500 ( .A0(n11322), .A1(n12763), .B0(n8393), .B1(n12762), .Y(
        n11321) );
  NOR2X1 U10501 ( .A(n8401), .B(n7976), .Y(n11322) );
  AOI22X1 U10502 ( .A0(n12751), .A1(n7879), .B0(n12755), .B1(test_se), .Y(
        n11320) );
  NAND2X1 U10503 ( .A(n11323), .B(n11324), .Y(n6131) );
  MX2X1 U10504 ( .A(n11325), .B(n11326), .S0(n11327), .Y(n11324) );
  NOR2X1 U10505 ( .A(n7400), .B(n11328), .Y(n11327) );
  NAND2X1 U10506 ( .A(n11293), .B(n7466), .Y(n11328) );
  NAND2X1 U10507 ( .A(g35), .B(n11329), .Y(n11326) );
  NAND2X1 U10508 ( .A(n7936), .B(n7391), .Y(n11325) );
  AOI22X1 U10509 ( .A0(n12761), .A1(n7879), .B0(n12763), .B1(test_se), .Y(
        n11323) );
  OAI21X1 U10510 ( .A0(n7866), .A1(n7347), .B0(n11330), .Y(n6130) );
  AOI22X1 U10511 ( .A0(n12753), .A1(n11331), .B0(n11314), .B1(n12754), .Y(
        n11330) );
  OAI21X1 U10512 ( .A0(n11332), .A1(n11333), .B0(n7920), .Y(n11331) );
  OAI21X1 U10513 ( .A0(n7921), .A1(n7210), .B0(n11334), .Y(n6129) );
  AOI21X1 U10514 ( .A0(n11314), .A1(n12752), .B0(n11335), .Y(n11334) );
  AOI21X1 U10515 ( .A0(n7866), .A1(n11336), .B0(n7550), .Y(n11335) );
  INVX1 U10516 ( .A(n11313), .Y(n11336) );
  NAND2X1 U10517 ( .A(n11337), .B(n11338), .Y(n6128) );
  MX2X1 U10518 ( .A(n7210), .B(n11305), .S0(n7852), .Y(n11338) );
  AOI22X1 U10519 ( .A0(n12764), .A1(n8393), .B0(n12762), .B1(n7879), .Y(n11337) );
  NOR2X1 U10520 ( .A(n11293), .B(n7976), .Y(n8393) );
  NAND2X1 U10521 ( .A(n11339), .B(n11340), .Y(n6127) );
  MX2X1 U10522 ( .A(n11341), .B(n11300), .S0(n11342), .Y(n11340) );
  NOR2X1 U10523 ( .A(n7400), .B(n11294), .Y(n11342) );
  NAND2X1 U10524 ( .A(n12764), .B(n11293), .Y(n11294) );
  NAND2X1 U10525 ( .A(n12757), .B(n7936), .Y(n11341) );
  AOI22X1 U10526 ( .A0(n12758), .A1(n7879), .B0(n12759), .B1(test_se), .Y(
        n11339) );
  NAND2X1 U10527 ( .A(n11343), .B(n11344), .Y(n6126) );
  MX2X1 U10528 ( .A(n11345), .B(n11300), .S0(n11346), .Y(n11344) );
  NOR2X1 U10529 ( .A(n12763), .B(n11305), .Y(n11346) );
  NAND2X1 U10530 ( .A(n12762), .B(n11293), .Y(n11305) );
  INVX1 U10531 ( .A(n8401), .Y(n11293) );
  NAND2X1 U10532 ( .A(n7936), .B(n11329), .Y(n11300) );
  NAND2X1 U10533 ( .A(n12893), .B(n8402), .Y(n11329) );
  NAND2X1 U10534 ( .A(n12758), .B(n7936), .Y(n11345) );
  AOI22X1 U10535 ( .A0(n7879), .A1(n7448), .B0(n12757), .B1(test_se), .Y(
        n11343) );
  NAND3X1 U10536 ( .A(n11347), .B(n11348), .C(n11349), .Y(n6125) );
  AOI22X1 U10537 ( .A0(n12752), .A1(n7879), .B0(n12764), .B1(test_se), .Y(
        n11349) );
  NAND2X1 U10538 ( .A(n11314), .B(n13022), .Y(n11348) );
  AOI22X1 U10539 ( .A0(n11350), .A1(n11351), .B0(n11313), .B1(n11352), .Y(
        n11347) );
  NAND3X1 U10540 ( .A(n11353), .B(n11354), .C(n11355), .Y(n11352) );
  AOI22X1 U10541 ( .A0(n11315), .A1(n7391), .B0(n11356), .B1(n12761), .Y(
        n11355) );
  NAND3X1 U10542 ( .A(n7485), .B(n7287), .C(n12757), .Y(n11354) );
  OR2X1 U10543 ( .A(n12754), .B(n11357), .Y(n11353) );
  AOI22X1 U10544 ( .A0(n12759), .A1(n12752), .B0(n12753), .B1(n12758), .Y(
        n11357) );
  INVX1 U10545 ( .A(n11319), .Y(n11351) );
  NAND3X1 U10546 ( .A(n12754), .B(n7287), .C(n11358), .Y(n11319) );
  NOR2X1 U10547 ( .A(n12756), .B(n7976), .Y(n11350) );
  NAND2X1 U10548 ( .A(n11359), .B(n11360), .Y(n6124) );
  MX2X1 U10549 ( .A(n11361), .B(n11362), .S0(n7594), .Y(n11360) );
  NAND2X1 U10550 ( .A(n11363), .B(n7936), .Y(n11362) );
  AOI21X1 U10551 ( .A0(n11364), .A1(n11365), .B0(n7879), .Y(n11361) );
  NOR2X1 U10552 ( .A(n11332), .B(n11363), .Y(n11364) );
  NOR2X1 U10553 ( .A(n12748), .B(n11315), .Y(n11363) );
  AOI22X1 U10554 ( .A0(n11314), .A1(n7436), .B0(n12760), .B1(test_se), .Y(
        n11359) );
  OAI21X1 U10555 ( .A0(n12748), .A1(n8721), .B0(n11366), .Y(n6123) );
  AOI22X1 U10556 ( .A0(n11367), .A1(n11368), .B0(n12747), .B1(n11369), .Y(
        n11366) );
  OAI21X1 U10557 ( .A0(n11315), .A1(n7976), .B0(n11370), .Y(n11369) );
  INVX1 U10558 ( .A(n11314), .Y(n11370) );
  XOR2X1 U10559 ( .A(n12760), .B(n7436), .Y(n11368) );
  AND2X1 U10560 ( .A(n11313), .B(n11315), .Y(n11367) );
  NOR2X1 U10561 ( .A(n7550), .B(n12753), .Y(n11315) );
  OAI21X1 U10562 ( .A0(n7936), .A1(n7351), .B0(n11371), .Y(n6122) );
  MX2X1 U10563 ( .A(n11372), .B(n11373), .S0(n7588), .Y(n11371) );
  NAND2X1 U10564 ( .A(n11356), .B(n11313), .Y(n11373) );
  MX2X1 U10565 ( .A(n12745), .B(n12746), .S0(n11295), .Y(n6121) );
  OAI21X1 U10566 ( .A0(n11295), .A1(n7237), .B0(n11374), .Y(n6120) );
  MX2X1 U10567 ( .A(n11375), .B(n11376), .S0(n12745), .Y(n11374) );
  AOI21X1 U10568 ( .A0(n12746), .A1(n8399), .B0(n8593), .Y(n11376) );
  NAND3X1 U10569 ( .A(n7936), .B(n7588), .C(n8399), .Y(n11375) );
  OAI21X1 U10570 ( .A0(n11295), .A1(n7309), .B0(n11377), .Y(n6119) );
  MX2X1 U10571 ( .A(n11378), .B(n7237), .S0(n7951), .Y(n11377) );
  NAND2X1 U10572 ( .A(n8399), .B(n7309), .Y(n11378) );
  INVX1 U10573 ( .A(n11299), .Y(n11295) );
  NOR2X1 U10574 ( .A(n7976), .B(n8399), .Y(n11299) );
  NOR2X1 U10575 ( .A(n8397), .B(n8401), .Y(n8399) );
  NOR2X1 U10576 ( .A(n11379), .B(n11380), .Y(n8401) );
  INVX1 U10577 ( .A(n8402), .Y(n11380) );
  NOR2X1 U10578 ( .A(n11282), .B(n12909), .Y(n8402) );
  AOI21X1 U10579 ( .A0(n11283), .A1(n10824), .B0(n7911), .Y(n11379) );
  NOR2X1 U10580 ( .A(n7551), .B(n12973), .Y(n10824) );
  OR2X1 U10581 ( .A(n12763), .B(n12764), .Y(n8397) );
  OAI22X1 U10582 ( .A0(n11372), .A1(n7663), .B0(n11381), .B1(n7309), .Y(n6118)
         );
  AOI21X1 U10583 ( .A0(n11356), .A1(n11358), .B0(n8593), .Y(n11381) );
  OAI21X1 U10584 ( .A0(n11372), .A1(n7212), .B0(n11382), .Y(n6117) );
  MX2X1 U10585 ( .A(n11383), .B(n11384), .S0(n7663), .Y(n11382) );
  NAND3X1 U10586 ( .A(n11313), .B(n7309), .C(n11356), .Y(n11384) );
  NOR2X1 U10587 ( .A(n11385), .B(n7976), .Y(n11313) );
  AOI21X1 U10588 ( .A0(n11386), .A1(n12744), .B0(n8593), .Y(n11383) );
  NOR2X1 U10589 ( .A(n11385), .B(n11387), .Y(n11386) );
  INVX1 U10590 ( .A(n11358), .Y(n11385) );
  AOI21X1 U10591 ( .A0(n11387), .A1(n7936), .B0(n11314), .Y(n11372) );
  NOR2X1 U10592 ( .A(n7976), .B(n11358), .Y(n11314) );
  NOR2X1 U10593 ( .A(n11388), .B(n11332), .Y(n11358) );
  AOI21X1 U10594 ( .A0(n11389), .A1(n13018), .B0(n11390), .Y(n11332) );
  INVX1 U10595 ( .A(n11356), .Y(n11387) );
  NOR2X1 U10596 ( .A(n7485), .B(n7287), .Y(n11356) );
  OAI22X1 U10597 ( .A0(n7866), .A1(n7212), .B0(n11391), .B1(n7976), .Y(n6116)
         );
  AOI22X1 U10598 ( .A0(n11392), .A1(n11393), .B0(n12742), .B1(n11394), .Y(
        n11391) );
  NOR2X1 U10599 ( .A(n12741), .B(n12743), .Y(n11392) );
  MX2X1 U10600 ( .A(n12739), .B(n12728), .S0(n11395), .Y(n6115) );
  NAND2X1 U10601 ( .A(n11396), .B(n11397), .Y(n6114) );
  AOI22X1 U10602 ( .A0(n11398), .A1(n8386), .B0(n12740), .B1(n11399), .Y(
        n11397) );
  INVX1 U10603 ( .A(n11400), .Y(n11398) );
  AOI22X1 U10604 ( .A0(n12739), .A1(n7879), .B0(test_se), .B1(n7392), .Y(
        n11396) );
  NAND2X1 U10605 ( .A(n11401), .B(n11402), .Y(n6113) );
  MX2X1 U10606 ( .A(n11403), .B(n11400), .S0(n11404), .Y(n11402) );
  NOR2X1 U10607 ( .A(n12743), .B(n11405), .Y(n11404) );
  NAND2X1 U10608 ( .A(n12738), .B(n7936), .Y(n11403) );
  AOI22X1 U10609 ( .A0(n7879), .A1(n7392), .B0(n12740), .B1(test_se), .Y(
        n11401) );
  NAND2X1 U10610 ( .A(n11406), .B(n11407), .Y(n6112) );
  MX2X1 U10611 ( .A(n11408), .B(n11400), .S0(n11409), .Y(n11407) );
  NOR2X1 U10612 ( .A(n12741), .B(n11394), .Y(n11409) );
  NAND2X1 U10613 ( .A(n7936), .B(n7449), .Y(n11408) );
  AOI22X1 U10614 ( .A0(n12738), .A1(n7879), .B0(n12737), .B1(test_se), .Y(
        n11406) );
  NAND2X1 U10615 ( .A(n11410), .B(n11411), .Y(n6111) );
  AOI22X1 U10616 ( .A0(n11412), .A1(n11413), .B0(n12732), .B1(n11414), .Y(
        n11411) );
  NOR2X1 U10617 ( .A(n12731), .B(n11415), .Y(n11412) );
  AOI22X1 U10618 ( .A0(n12734), .A1(n7879), .B0(test_se), .B1(n7449), .Y(
        n11410) );
  OAI21X1 U10619 ( .A0(n7866), .A1(n7486), .B0(n11416), .Y(n6110) );
  AOI22X1 U10620 ( .A0(n11417), .A1(n7936), .B0(n12736), .B1(n7879), .Y(n11416) );
  MX2X1 U10621 ( .A(n11418), .B(n12734), .S0(n11419), .Y(n11417) );
  NAND2X1 U10622 ( .A(n12741), .B(n7401), .Y(n11418) );
  NAND2X1 U10623 ( .A(n11420), .B(n11421), .Y(n6109) );
  AOI22X1 U10624 ( .A0(n11422), .A1(n12742), .B0(n8380), .B1(n12741), .Y(
        n11421) );
  NOR2X1 U10625 ( .A(n8388), .B(n7976), .Y(n11422) );
  AOI22X1 U10626 ( .A0(n12730), .A1(n7878), .B0(n12734), .B1(test_se), .Y(
        n11420) );
  NAND2X1 U10627 ( .A(n11423), .B(n11424), .Y(n6108) );
  MX2X1 U10628 ( .A(n11425), .B(n11426), .S0(n11427), .Y(n11424) );
  NOR2X1 U10629 ( .A(n7401), .B(n11428), .Y(n11427) );
  NAND2X1 U10630 ( .A(n11393), .B(n7467), .Y(n11428) );
  NAND2X1 U10631 ( .A(g35), .B(n11429), .Y(n11426) );
  NAND2X1 U10632 ( .A(n7936), .B(n7392), .Y(n11425) );
  AOI22X1 U10633 ( .A0(n12740), .A1(n7878), .B0(n12742), .B1(test_se), .Y(
        n11423) );
  OAI21X1 U10634 ( .A0(n7865), .A1(n7694), .B0(n11430), .Y(n6107) );
  AOI22X1 U10635 ( .A0(n12732), .A1(n11431), .B0(n11414), .B1(n12733), .Y(
        n11430) );
  OAI21X1 U10636 ( .A0(n11432), .A1(n11433), .B0(n7920), .Y(n11431) );
  OAI21X1 U10637 ( .A0(n7865), .A1(n7288), .B0(n11434), .Y(n6106) );
  AOI22X1 U10638 ( .A0(n12733), .A1(n7878), .B0(n12729), .B1(n7936), .Y(n11434) );
  OAI21X1 U10639 ( .A0(n7921), .A1(n7235), .B0(n11435), .Y(n6105) );
  AOI21X1 U10640 ( .A0(n12731), .A1(n11414), .B0(n11436), .Y(n11435) );
  AOI21X1 U10641 ( .A0(n7865), .A1(n11437), .B0(n7552), .Y(n11436) );
  INVX1 U10642 ( .A(n11413), .Y(n11437) );
  NAND2X1 U10643 ( .A(n11438), .B(n11439), .Y(n6104) );
  MX2X1 U10644 ( .A(n7235), .B(n11405), .S0(n7852), .Y(n11439) );
  AOI22X1 U10645 ( .A0(n12743), .A1(n8380), .B0(n12741), .B1(n7878), .Y(n11438) );
  NOR2X1 U10646 ( .A(n11393), .B(n7974), .Y(n8380) );
  NAND2X1 U10647 ( .A(n11440), .B(n11441), .Y(n6103) );
  MX2X1 U10648 ( .A(n11442), .B(n11400), .S0(n11443), .Y(n11441) );
  NOR2X1 U10649 ( .A(n7401), .B(n11394), .Y(n11443) );
  NAND2X1 U10650 ( .A(n12743), .B(n11393), .Y(n11394) );
  NAND2X1 U10651 ( .A(n12736), .B(n7936), .Y(n11442) );
  AOI22X1 U10652 ( .A0(n12737), .A1(n7878), .B0(n12738), .B1(test_se), .Y(
        n11440) );
  NAND2X1 U10653 ( .A(n11444), .B(n11445), .Y(n6102) );
  MX2X1 U10654 ( .A(n11446), .B(n11400), .S0(n11447), .Y(n11445) );
  NOR2X1 U10655 ( .A(n12742), .B(n11405), .Y(n11447) );
  NAND2X1 U10656 ( .A(n12741), .B(n11393), .Y(n11405) );
  INVX1 U10657 ( .A(n8388), .Y(n11393) );
  NAND2X1 U10658 ( .A(n7936), .B(n11429), .Y(n11400) );
  NAND2X1 U10659 ( .A(n8389), .B(n7474), .Y(n11429) );
  NAND2X1 U10660 ( .A(n12737), .B(n7936), .Y(n11446) );
  AOI22X1 U10661 ( .A0(n7878), .A1(n7449), .B0(n12736), .B1(test_se), .Y(
        n11444) );
  NAND3X1 U10662 ( .A(n11448), .B(n11449), .C(n11450), .Y(n6101) );
  AOI22X1 U10663 ( .A0(n12731), .A1(n7878), .B0(n12743), .B1(test_se), .Y(
        n11450) );
  NAND2X1 U10664 ( .A(n11414), .B(n13024), .Y(n11449) );
  AOI22X1 U10665 ( .A0(n11451), .A1(n11452), .B0(n11413), .B1(n11453), .Y(
        n11448) );
  NAND3X1 U10666 ( .A(n11454), .B(n11455), .C(n11456), .Y(n11453) );
  AOI22X1 U10667 ( .A0(n11415), .A1(n7392), .B0(n11457), .B1(n12740), .Y(
        n11456) );
  NAND3X1 U10668 ( .A(n7486), .B(n7288), .C(n12736), .Y(n11455) );
  OR2X1 U10669 ( .A(n12733), .B(n11458), .Y(n11454) );
  AOI22X1 U10670 ( .A0(n12731), .A1(n12738), .B0(n12732), .B1(n12737), .Y(
        n11458) );
  INVX1 U10671 ( .A(n11419), .Y(n11452) );
  NAND3X1 U10672 ( .A(n11459), .B(n7288), .C(n12733), .Y(n11419) );
  NOR2X1 U10673 ( .A(n12735), .B(n7974), .Y(n11451) );
  NAND2X1 U10674 ( .A(n11460), .B(n11461), .Y(n6100) );
  MX2X1 U10675 ( .A(n11462), .B(n11463), .S0(n7595), .Y(n11461) );
  NAND2X1 U10676 ( .A(n11464), .B(n7936), .Y(n11463) );
  AOI21X1 U10677 ( .A0(n11465), .A1(n11466), .B0(n7878), .Y(n11462) );
  NOR2X1 U10678 ( .A(n11432), .B(n11464), .Y(n11465) );
  NOR2X1 U10679 ( .A(n12727), .B(n11415), .Y(n11464) );
  AOI22X1 U10680 ( .A0(n11414), .A1(n7437), .B0(n12739), .B1(test_se), .Y(
        n11460) );
  OAI21X1 U10681 ( .A0(n12727), .A1(n8721), .B0(n11467), .Y(n6099) );
  AOI22X1 U10682 ( .A0(n11468), .A1(n11469), .B0(n12726), .B1(n11470), .Y(
        n11467) );
  OAI21X1 U10683 ( .A0(n11415), .A1(n7974), .B0(n11471), .Y(n11470) );
  INVX1 U10684 ( .A(n11414), .Y(n11471) );
  XOR2X1 U10685 ( .A(n12739), .B(n7437), .Y(n11469) );
  AND2X1 U10686 ( .A(n11413), .B(n11415), .Y(n11468) );
  NOR2X1 U10687 ( .A(n7552), .B(n12732), .Y(n11415) );
  OAI21X1 U10688 ( .A0(n7936), .A1(n7241), .B0(n11472), .Y(n6098) );
  MX2X1 U10689 ( .A(n11473), .B(n11474), .S0(n7589), .Y(n11472) );
  NAND2X1 U10690 ( .A(n11457), .B(n11413), .Y(n11474) );
  MX2X1 U10691 ( .A(n12724), .B(n12725), .S0(n11395), .Y(n6097) );
  OAI21X1 U10692 ( .A0(n11395), .A1(n7648), .B0(n11475), .Y(n6096) );
  MX2X1 U10693 ( .A(n11476), .B(n11477), .S0(n12724), .Y(n11475) );
  AOI21X1 U10694 ( .A0(n12725), .A1(n8386), .B0(n8593), .Y(n11477) );
  NAND3X1 U10695 ( .A(n7936), .B(n7589), .C(n8386), .Y(n11476) );
  OAI21X1 U10696 ( .A0(n11395), .A1(n7310), .B0(n11478), .Y(n6095) );
  MX2X1 U10697 ( .A(n11479), .B(n7648), .S0(n7955), .Y(n11478) );
  NAND2X1 U10698 ( .A(n8386), .B(n7310), .Y(n11479) );
  INVX1 U10699 ( .A(n11399), .Y(n11395) );
  NOR2X1 U10700 ( .A(n7974), .B(n8386), .Y(n11399) );
  NOR2X1 U10701 ( .A(n8384), .B(n8388), .Y(n8386) );
  NOR2X1 U10702 ( .A(n11480), .B(n11481), .Y(n8388) );
  INVX1 U10703 ( .A(n8389), .Y(n11481) );
  NOR2X1 U10704 ( .A(n11282), .B(n12908), .Y(n8389) );
  AOI21X1 U10705 ( .A0(n10719), .A1(n11283), .B0(n699), .Y(n11480) );
  INVX1 U10706 ( .A(n10718), .Y(n10719) );
  NAND2X1 U10707 ( .A(n12973), .B(n12972), .Y(n10718) );
  OR2X1 U10708 ( .A(n12742), .B(n12743), .Y(n8384) );
  OAI22X1 U10709 ( .A0(n11473), .A1(n7664), .B0(n11482), .B1(n7310), .Y(n6094)
         );
  AOI21X1 U10710 ( .A0(n11457), .A1(n11459), .B0(n8593), .Y(n11482) );
  OAI21X1 U10711 ( .A0(n11473), .A1(n7336), .B0(n11483), .Y(n6093) );
  MX2X1 U10712 ( .A(n11484), .B(n11485), .S0(n7664), .Y(n11483) );
  NAND3X1 U10713 ( .A(n11413), .B(n7310), .C(n11457), .Y(n11485) );
  NOR2X1 U10714 ( .A(n11486), .B(n7974), .Y(n11413) );
  AOI21X1 U10715 ( .A0(n11487), .A1(n12723), .B0(n8593), .Y(n11484) );
  NOR2X1 U10716 ( .A(n11486), .B(n11488), .Y(n11487) );
  INVX1 U10717 ( .A(n11459), .Y(n11486) );
  AOI21X1 U10718 ( .A0(n11488), .A1(n7936), .B0(n11414), .Y(n11473) );
  NOR2X1 U10719 ( .A(n7974), .B(n11459), .Y(n11414) );
  NOR2X1 U10720 ( .A(n11489), .B(n11432), .Y(n11459) );
  AOI21X1 U10721 ( .A0(n11389), .A1(n13021), .B0(n11390), .Y(n11432) );
  INVX1 U10722 ( .A(n11457), .Y(n11488) );
  NOR2X1 U10723 ( .A(n7288), .B(n7486), .Y(n11457) );
  OAI22X1 U10724 ( .A0(n7865), .A1(n7336), .B0(n11490), .B1(n7974), .Y(n6092)
         );
  AOI22X1 U10725 ( .A0(n11491), .A1(n11492), .B0(n12721), .B1(n11493), .Y(
        n11490) );
  NOR2X1 U10726 ( .A(n12720), .B(n12722), .Y(n11491) );
  MX2X1 U10727 ( .A(n12718), .B(n12707), .S0(n11208), .Y(n6091) );
  INVX1 U10728 ( .A(n11494), .Y(n11208) );
  NAND2X1 U10729 ( .A(n11495), .B(n11496), .Y(n6090) );
  AOI22X1 U10730 ( .A0(n11494), .A1(n12719), .B0(n11497), .B1(n8373), .Y(
        n11496) );
  INVX1 U10731 ( .A(n11498), .Y(n11497) );
  NOR2X1 U10732 ( .A(n7974), .B(n8373), .Y(n11494) );
  NOR2X1 U10733 ( .A(n8371), .B(n8375), .Y(n8373) );
  OR2X1 U10734 ( .A(n12721), .B(n12722), .Y(n8371) );
  AOI22X1 U10735 ( .A0(n12718), .A1(n7878), .B0(test_se), .B1(n7393), .Y(
        n11495) );
  NAND2X1 U10736 ( .A(n11499), .B(n11500), .Y(n6089) );
  MX2X1 U10737 ( .A(n11501), .B(n11498), .S0(n11502), .Y(n11500) );
  NOR2X1 U10738 ( .A(n12722), .B(n11503), .Y(n11502) );
  NAND2X1 U10739 ( .A(n12717), .B(n7936), .Y(n11501) );
  AOI22X1 U10740 ( .A0(n7878), .A1(n7393), .B0(n12719), .B1(test_se), .Y(
        n11499) );
  NAND2X1 U10741 ( .A(n11504), .B(n11505), .Y(n6088) );
  MX2X1 U10742 ( .A(n11506), .B(n11498), .S0(n11507), .Y(n11505) );
  NOR2X1 U10743 ( .A(n12720), .B(n11493), .Y(n11507) );
  NAND2X1 U10744 ( .A(n7936), .B(n7450), .Y(n11506) );
  AOI22X1 U10745 ( .A0(n12717), .A1(n7878), .B0(n12716), .B1(test_se), .Y(
        n11504) );
  NAND2X1 U10746 ( .A(n11508), .B(n11509), .Y(n6087) );
  MX2X1 U10747 ( .A(n11510), .B(n11498), .S0(n11511), .Y(n11509) );
  NOR2X1 U10748 ( .A(n12721), .B(n11503), .Y(n11511) );
  NAND2X1 U10749 ( .A(n12716), .B(n7936), .Y(n11510) );
  AOI22X1 U10750 ( .A0(n7878), .A1(n7450), .B0(n12715), .B1(test_se), .Y(
        n11508) );
  NAND2X1 U10751 ( .A(n11512), .B(n11513), .Y(n6086) );
  MX2X1 U10752 ( .A(n11514), .B(n11498), .S0(n11515), .Y(n11513) );
  NOR2X1 U10753 ( .A(n7402), .B(n11493), .Y(n11515) );
  NAND2X1 U10754 ( .A(n12722), .B(n11492), .Y(n11493) );
  NAND2X1 U10755 ( .A(n7937), .B(n11516), .Y(n11498) );
  NAND2X1 U10756 ( .A(n12715), .B(n7937), .Y(n11514) );
  AOI22X1 U10757 ( .A0(n12716), .A1(n7876), .B0(n12717), .B1(test_se), .Y(
        n11512) );
  OAI21X1 U10758 ( .A0(n7865), .A1(n7487), .B0(n11517), .Y(n6085) );
  AOI22X1 U10759 ( .A0(n11518), .A1(n7937), .B0(n12715), .B1(n7876), .Y(n11517) );
  MX2X1 U10760 ( .A(n11519), .B(n12713), .S0(n11192), .Y(n11518) );
  NAND3X1 U10761 ( .A(n11215), .B(n7289), .C(n12712), .Y(n11192) );
  NAND2X1 U10762 ( .A(n12720), .B(n7402), .Y(n11519) );
  NAND2X1 U10763 ( .A(n11520), .B(n11521), .Y(n6084) );
  AOI22X1 U10764 ( .A0(n11522), .A1(n12721), .B0(n8367), .B1(n12720), .Y(
        n11521) );
  NOR2X1 U10765 ( .A(n8375), .B(n7974), .Y(n11522) );
  AOI22X1 U10766 ( .A0(n12709), .A1(n7876), .B0(n12713), .B1(test_se), .Y(
        n11520) );
  NAND2X1 U10767 ( .A(n11523), .B(n11524), .Y(n6083) );
  MX2X1 U10768 ( .A(n11525), .B(n11526), .S0(n11527), .Y(n11524) );
  NOR2X1 U10769 ( .A(n7402), .B(n11528), .Y(n11527) );
  NAND2X1 U10770 ( .A(n11492), .B(n7468), .Y(n11528) );
  NAND2X1 U10771 ( .A(g35), .B(n11516), .Y(n11526) );
  OR2X1 U10772 ( .A(n7474), .B(n8376), .Y(n11516) );
  NAND2X1 U10773 ( .A(n7937), .B(n7393), .Y(n11525) );
  AOI22X1 U10774 ( .A0(n12719), .A1(n7876), .B0(n12721), .B1(test_se), .Y(
        n11523) );
  OAI21X1 U10775 ( .A0(n7865), .A1(n7348), .B0(n11529), .Y(n6082) );
  AOI22X1 U10776 ( .A0(n12711), .A1(n11530), .B0(n11179), .B1(n12712), .Y(
        n11529) );
  OAI21X1 U10777 ( .A0(n11199), .A1(n11531), .B0(n7920), .Y(n11530) );
  OAI21X1 U10778 ( .A0(n7865), .A1(n7289), .B0(n11532), .Y(n6081) );
  AOI22X1 U10779 ( .A0(n12712), .A1(n7876), .B0(n12708), .B1(n7937), .Y(n11532) );
  OAI21X1 U10780 ( .A0(n7921), .A1(n7211), .B0(n11533), .Y(n6080) );
  AOI21X1 U10781 ( .A0(n12710), .A1(n11179), .B0(n11534), .Y(n11533) );
  AOI21X1 U10782 ( .A0(n7865), .A1(n11535), .B0(n7553), .Y(n11534) );
  INVX1 U10783 ( .A(n11178), .Y(n11535) );
  NOR2X1 U10784 ( .A(n11220), .B(n7974), .Y(n11178) );
  INVX1 U10785 ( .A(n11215), .Y(n11220) );
  NOR2X1 U10786 ( .A(n7974), .B(n11215), .Y(n11179) );
  NOR2X1 U10787 ( .A(n11536), .B(n11199), .Y(n11215) );
  AOI21X1 U10788 ( .A0(n11389), .A1(n13019), .B0(n11390), .Y(n11199) );
  NAND2X1 U10789 ( .A(n11537), .B(n11538), .Y(n6079) );
  MX2X1 U10790 ( .A(n7211), .B(n11503), .S0(n7852), .Y(n11538) );
  NAND2X1 U10791 ( .A(n12720), .B(n11492), .Y(n11503) );
  AOI22X1 U10792 ( .A0(n12722), .A1(n8367), .B0(n12720), .B1(n7876), .Y(n11537) );
  NOR2X1 U10793 ( .A(n11492), .B(n7974), .Y(n8367) );
  INVX1 U10794 ( .A(n8375), .Y(n11492) );
  NOR2X1 U10795 ( .A(n11539), .B(n8376), .Y(n8375) );
  OR2X1 U10796 ( .A(n11282), .B(n12968), .Y(n8376) );
  NAND2X1 U10797 ( .A(n8779), .B(n8783), .Y(n11282) );
  AOI21X1 U10798 ( .A0(n11283), .A1(n10713), .B0(n7313), .Y(n11539) );
  NOR2X1 U10799 ( .A(n12972), .B(n12973), .Y(n10713) );
  INVX1 U10800 ( .A(n11540), .Y(n11283) );
  NAND4X1 U10801 ( .A(n11541), .B(n12941), .C(n11542), .D(n7509), .Y(n11540)
         );
  NOR2X1 U10802 ( .A(n12897), .B(n12942), .Y(n11542) );
  NOR2X1 U10803 ( .A(n7256), .B(n7479), .Y(n11541) );
  NAND3X1 U10804 ( .A(n11543), .B(n11544), .C(n11545), .Y(n6078) );
  AOI22X1 U10805 ( .A0(n12780), .A1(n7876), .B0(n12793), .B1(test_se), .Y(
        n11545) );
  NAND2X1 U10806 ( .A(n8760), .B(n13025), .Y(n11544) );
  NOR2X1 U10807 ( .A(n7974), .B(n8758), .Y(n8760) );
  AOI22X1 U10808 ( .A0(n11546), .A1(n11547), .B0(n8766), .B1(n11548), .Y(
        n11543) );
  NAND3X1 U10809 ( .A(n11549), .B(n11550), .C(n11551), .Y(n11548) );
  AOI22X1 U10810 ( .A0(n12790), .A1(n8759), .B0(n11274), .B1(n12789), .Y(
        n11551) );
  NOR2X1 U10811 ( .A(n7457), .B(n7290), .Y(n11274) );
  NOR2X1 U10812 ( .A(n7488), .B(n12782), .Y(n8759) );
  NAND3X1 U10813 ( .A(n7457), .B(n7290), .C(n12785), .Y(n11550) );
  OR2X1 U10814 ( .A(n12781), .B(n11552), .Y(n11549) );
  AOI22X1 U10815 ( .A0(n12787), .A1(n12780), .B0(n12786), .B1(n12782), .Y(
        n11552) );
  NOR2X1 U10816 ( .A(n11231), .B(n7972), .Y(n8766) );
  INVX1 U10817 ( .A(n8758), .Y(n11231) );
  INVX1 U10818 ( .A(n11225), .Y(n11547) );
  NAND3X1 U10819 ( .A(n12781), .B(n7290), .C(n8758), .Y(n11225) );
  NOR2X1 U10820 ( .A(n11553), .B(n11554), .Y(n8758) );
  AOI21X1 U10821 ( .A0(n13020), .A1(n11389), .B0(n11390), .Y(n11553) );
  NOR2X1 U10822 ( .A(n12784), .B(n7972), .Y(n11546) );
  OR2X1 U10823 ( .A(n13030), .B(n7937), .Y(n6077) );
  OAI21X1 U10824 ( .A0(n13011), .A1(n7865), .B0(n11555), .Y(n6076) );
  AOI22X1 U10825 ( .A0(n11556), .A1(n7937), .B0(n12698), .B1(n7876), .Y(n11555) );
  INVX1 U10826 ( .A(n11557), .Y(n11556) );
  MX2X1 U10827 ( .A(n7531), .B(n12698), .S0(n11174), .Y(n11557) );
  AND2X1 U10828 ( .A(n11558), .B(n11559), .Y(n11174) );
  NAND2X1 U10829 ( .A(n11560), .B(n11561), .Y(n6075) );
  AOI22X1 U10830 ( .A0(n11562), .A1(n8732), .B0(n12804), .B1(n8720), .Y(n11561) );
  NOR2X1 U10831 ( .A(n12802), .B(n8719), .Y(n11562) );
  AOI22X1 U10832 ( .A0(n12805), .A1(n7876), .B0(test_se), .B1(n7451), .Y(
        n11560) );
  OAI21X1 U10833 ( .A0(n7865), .A1(n7489), .B0(n11563), .Y(n6074) );
  AOI22X1 U10834 ( .A0(n11564), .A1(n7937), .B0(n12807), .B1(n7876), .Y(n11563) );
  MX2X1 U10835 ( .A(n11565), .B(n12805), .S0(n11566), .Y(n11564) );
  NAND2X1 U10836 ( .A(n12818), .B(n7403), .Y(n11565) );
  OAI21X1 U10837 ( .A0(n7865), .A1(n7687), .B0(n11567), .Y(n6073) );
  AOI22X1 U10838 ( .A0(n11568), .A1(n7937), .B0(n12801), .B1(n7876), .Y(n11567) );
  MX2X1 U10839 ( .A(n12818), .B(n12819), .S0(n8708), .Y(n11568) );
  OAI21X1 U10840 ( .A0(n7865), .A1(n7469), .B0(n11569), .Y(n6072) );
  AOI22X1 U10841 ( .A0(n12819), .A1(n7876), .B0(n12801), .B1(n7937), .Y(n11569) );
  OAI21X1 U10842 ( .A0(n7865), .A1(n7346), .B0(n11570), .Y(n6071) );
  AOI22X1 U10843 ( .A0(n12804), .A1(n11571), .B0(n12803), .B1(n8720), .Y(
        n11570) );
  OAI21X1 U10844 ( .A0(n8718), .A1(n11531), .B0(n7920), .Y(n11571) );
  INVX1 U10845 ( .A(n8717), .Y(n11531) );
  NOR2X1 U10846 ( .A(n11536), .B(test_se), .Y(n8717) );
  OAI21X1 U10847 ( .A0(n7865), .A1(n7291), .B0(n11572), .Y(n6070) );
  AOI22X1 U10848 ( .A0(n12803), .A1(n7875), .B0(n12800), .B1(n7937), .Y(n11572) );
  OAI21X1 U10849 ( .A0(n7921), .A1(n7209), .B0(n11573), .Y(n6069) );
  AOI21X1 U10850 ( .A0(n12802), .A1(n8720), .B0(n11574), .Y(n11573) );
  AOI21X1 U10851 ( .A0(n7865), .A1(n8727), .B0(n7554), .Y(n11574) );
  INVX1 U10852 ( .A(n8732), .Y(n8727) );
  NAND2X1 U10853 ( .A(n11575), .B(n11576), .Y(n6068) );
  MX2X1 U10854 ( .A(n7209), .B(n11577), .S0(n7853), .Y(n11576) );
  AOI22X1 U10855 ( .A0(n11578), .A1(n8423), .B0(n12818), .B1(n7875), .Y(n11575) );
  AND2X1 U10856 ( .A(n7937), .B(n12820), .Y(n11578) );
  NAND2X1 U10857 ( .A(n11579), .B(n11580), .Y(n6067) );
  AOI22X1 U10858 ( .A0(n12811), .A1(n8738), .B0(n11581), .B1(n8424), .Y(n11580) );
  INVX1 U10859 ( .A(n11582), .Y(n11581) );
  NOR2X1 U10860 ( .A(n7972), .B(n8424), .Y(n8738) );
  NOR2X1 U10861 ( .A(n8422), .B(n8423), .Y(n8424) );
  INVX1 U10862 ( .A(n8708), .Y(n8423) );
  OR2X1 U10863 ( .A(n12819), .B(n12820), .Y(n8422) );
  AOI22X1 U10864 ( .A0(n12810), .A1(n7875), .B0(test_se), .B1(n7394), .Y(
        n11579) );
  NAND2X1 U10865 ( .A(n11583), .B(n11584), .Y(n6066) );
  MX2X1 U10866 ( .A(n11585), .B(n11586), .S0(n11587), .Y(n11584) );
  NOR2X1 U10867 ( .A(n7403), .B(n11588), .Y(n11587) );
  NAND2X1 U10868 ( .A(n8708), .B(n7469), .Y(n11588) );
  OAI21X1 U10869 ( .A0(n7362), .A1(n11589), .B0(g35), .Y(n11586) );
  NAND2X1 U10870 ( .A(n7937), .B(n7394), .Y(n11585) );
  AOI22X1 U10871 ( .A0(n12811), .A1(n7875), .B0(n12819), .B1(test_se), .Y(
        n11583) );
  NAND2X1 U10872 ( .A(n11590), .B(n11591), .Y(n6065) );
  MX2X1 U10873 ( .A(n11592), .B(n11582), .S0(n11593), .Y(n11591) );
  NOR2X1 U10874 ( .A(n12820), .B(n11577), .Y(n11593) );
  NAND2X1 U10875 ( .A(n12809), .B(n7937), .Y(n11592) );
  AOI22X1 U10876 ( .A0(n7875), .A1(n7394), .B0(n12811), .B1(test_se), .Y(
        n11590) );
  NAND2X1 U10877 ( .A(n11594), .B(n11595), .Y(n6064) );
  MX2X1 U10878 ( .A(n11596), .B(n11582), .S0(n11597), .Y(n11595) );
  NOR2X1 U10879 ( .A(n12818), .B(n8709), .Y(n11597) );
  NAND2X1 U10880 ( .A(n7937), .B(n7451), .Y(n11596) );
  AOI22X1 U10881 ( .A0(n12809), .A1(n7875), .B0(n12808), .B1(test_se), .Y(
        n11594) );
  NAND2X1 U10882 ( .A(n11598), .B(n11599), .Y(n6063) );
  MX2X1 U10883 ( .A(n11600), .B(n11582), .S0(n11601), .Y(n11599) );
  NOR2X1 U10884 ( .A(n12819), .B(n11577), .Y(n11601) );
  NAND2X1 U10885 ( .A(n12818), .B(n8708), .Y(n11577) );
  NAND2X1 U10886 ( .A(n12808), .B(n7937), .Y(n11600) );
  AOI22X1 U10887 ( .A0(n7875), .A1(n7451), .B0(n12807), .B1(test_se), .Y(
        n11598) );
  NAND2X1 U10888 ( .A(n11602), .B(n11603), .Y(n6062) );
  MX2X1 U10889 ( .A(n11604), .B(n11582), .S0(n11605), .Y(n11603) );
  NOR2X1 U10890 ( .A(n7403), .B(n8709), .Y(n11605) );
  NAND2X1 U10891 ( .A(n12820), .B(n8708), .Y(n8709) );
  NAND3X1 U10892 ( .A(n8452), .B(n11606), .C(n13035), .Y(n8708) );
  OAI21X1 U10893 ( .A0(n10626), .A1(n11607), .B0(n13048), .Y(n11606) );
  OR2X1 U10894 ( .A(n13053), .B(n13054), .Y(n10626) );
  OAI21X1 U10895 ( .A0(n7362), .A1(n11589), .B0(n7922), .Y(n11582) );
  NAND2X1 U10896 ( .A(n12807), .B(n7937), .Y(n11604) );
  AOI22X1 U10897 ( .A0(n12808), .A1(n7875), .B0(n12809), .B1(test_se), .Y(
        n11602) );
  NAND3X1 U10898 ( .A(n11608), .B(n11609), .C(n11610), .Y(n6061) );
  AOI22X1 U10899 ( .A0(n12802), .A1(n7875), .B0(n12820), .B1(test_se), .Y(
        n11610) );
  NAND2X1 U10900 ( .A(n8720), .B(n13013), .Y(n11609) );
  NOR2X1 U10901 ( .A(n7972), .B(n8740), .Y(n8720) );
  AOI22X1 U10902 ( .A0(n11611), .A1(n11612), .B0(n8732), .B1(n11613), .Y(
        n11608) );
  NAND3X1 U10903 ( .A(n11614), .B(n11615), .C(n11616), .Y(n11613) );
  AOI22X1 U10904 ( .A0(n8719), .A1(n7394), .B0(n12811), .B1(n8731), .Y(n11616)
         );
  NOR2X1 U10905 ( .A(n7291), .B(n7489), .Y(n8731) );
  NOR2X1 U10906 ( .A(n7554), .B(n12804), .Y(n8719) );
  NAND3X1 U10907 ( .A(n7489), .B(n7291), .C(n12807), .Y(n11615) );
  OR2X1 U10908 ( .A(n12803), .B(n11617), .Y(n11614) );
  AOI22X1 U10909 ( .A0(n12809), .A1(n12802), .B0(n12808), .B1(n12804), .Y(
        n11617) );
  NOR2X1 U10910 ( .A(n8745), .B(n7972), .Y(n8732) );
  INVX1 U10911 ( .A(n8740), .Y(n8745) );
  INVX1 U10912 ( .A(n11566), .Y(n11612) );
  NAND3X1 U10913 ( .A(n12803), .B(n7291), .C(n8740), .Y(n11566) );
  NOR2X1 U10914 ( .A(n11536), .B(n8718), .Y(n8740) );
  AOI21X1 U10915 ( .A0(n7531), .A1(n11389), .B0(n11390), .Y(n8718) );
  INVX1 U10916 ( .A(n11618), .Y(n11536) );
  NOR2X1 U10917 ( .A(n12806), .B(n7972), .Y(n11611) );
  NAND2X1 U10918 ( .A(n11619), .B(n11620), .Y(n6060) );
  AOI22X1 U10919 ( .A0(n11159), .A1(n7732), .B0(n11160), .B1(n7328), .Y(n11620) );
  AOI22X1 U10920 ( .A0(n7875), .A1(n7303), .B0(n13009), .B1(test_se), .Y(
        n11619) );
  OAI21X1 U10921 ( .A0(n12700), .A1(n7865), .B0(n11621), .Y(n6059) );
  AOI22X1 U10922 ( .A0(n11622), .A1(n7937), .B0(n13009), .B1(n7875), .Y(n11621) );
  MX2X1 U10923 ( .A(n7414), .B(n12699), .S0(n11171), .Y(n11622) );
  AND2X1 U10924 ( .A(n11623), .B(n11559), .Y(n11171) );
  OAI21X1 U10925 ( .A0(n13010), .A1(n7865), .B0(n11624), .Y(n6058) );
  AOI22X1 U10926 ( .A0(n11625), .A1(n7937), .B0(n7875), .B1(n7414), .Y(n11624)
         );
  MX2X1 U10927 ( .A(n12700), .B(n7377), .S0(n11166), .Y(n11625) );
  NAND3X1 U10928 ( .A(n11559), .B(n7300), .C(n13028), .Y(n11166) );
  INVX1 U10929 ( .A(n11626), .Y(n11559) );
  OAI21X1 U10930 ( .A0(n12701), .A1(n7865), .B0(n11627), .Y(n6057) );
  AOI22X1 U10931 ( .A0(n11628), .A1(n7937), .B0(n7905), .B1(n7377), .Y(n11627)
         );
  MX2X1 U10932 ( .A(n7297), .B(n12701), .S0(n11163), .Y(n11628) );
  NOR2X1 U10933 ( .A(n11626), .B(n11390), .Y(n11163) );
  NAND4X1 U10934 ( .A(n11629), .B(n11630), .C(n11631), .D(n11632), .Y(n6056)
         );
  OR2X1 U10935 ( .A(n11633), .B(n11634), .Y(n11632) );
  AOI21X1 U10936 ( .A0(n12887), .A1(n11635), .B0(n11636), .Y(n11633) );
  OAI21X1 U10937 ( .A0(n12879), .A1(n11637), .B0(n11638), .Y(n11636) );
  NAND3X1 U10938 ( .A(n7273), .B(n7404), .C(n12883), .Y(n11638) );
  AOI22X1 U10939 ( .A0(n12885), .A1(n12878), .B0(n12880), .B1(n12884), .Y(
        n11637) );
  AOI22X1 U10940 ( .A0(n11639), .A1(n11640), .B0(n11641), .B1(n11642), .Y(
        n11631) );
  NOR2X1 U10941 ( .A(n12882), .B(n7972), .Y(n11639) );
  NAND2X1 U10942 ( .A(n12890), .B(test_se), .Y(n11630) );
  AOI22X1 U10943 ( .A0(n11643), .A1(n13015), .B0(n12878), .B1(n7899), .Y(
        n11629) );
  MX2X1 U10944 ( .A(n12886), .B(n12875), .S0(n11644), .Y(n6055) );
  NAND2X1 U10945 ( .A(n11645), .B(n11646), .Y(n6054) );
  AOI22X1 U10946 ( .A0(n11647), .A1(n8461), .B0(n11648), .B1(n12887), .Y(
        n11646) );
  AOI22X1 U10947 ( .A0(n12886), .A1(n7900), .B0(n12888), .B1(test_se), .Y(
        n11645) );
  NAND2X1 U10948 ( .A(n11649), .B(n11650), .Y(n6053) );
  MX2X1 U10949 ( .A(n11651), .B(n11652), .S0(n11653), .Y(n11650) );
  NOR2X1 U10950 ( .A(n12890), .B(n11654), .Y(n11653) );
  NAND2X1 U10951 ( .A(n12885), .B(n7937), .Y(n11651) );
  AOI22X1 U10952 ( .A0(n12888), .A1(n7880), .B0(n12887), .B1(test_se), .Y(
        n11649) );
  NAND2X1 U10953 ( .A(n11655), .B(n11656), .Y(n6052) );
  MX2X1 U10954 ( .A(n11657), .B(n11652), .S0(n11658), .Y(n11656) );
  NOR2X1 U10955 ( .A(n11659), .B(n11660), .Y(n11658) );
  NAND2X1 U10956 ( .A(n7937), .B(n7452), .Y(n11657) );
  AOI22X1 U10957 ( .A0(n12885), .A1(n7906), .B0(n12884), .B1(test_se), .Y(
        n11655) );
  NAND2X1 U10958 ( .A(n11661), .B(n11662), .Y(n6051) );
  AOI22X1 U10959 ( .A0(n11663), .A1(n11664), .B0(n12880), .B1(n11665), .Y(
        n11662) );
  NOR2X1 U10960 ( .A(n12878), .B(n12879), .Y(n11663) );
  AOI22X1 U10961 ( .A0(n12881), .A1(n7898), .B0(test_se), .B1(n7452), .Y(
        n11661) );
  OAI21X1 U10962 ( .A0(n7865), .A1(n7273), .B0(n11666), .Y(n6050) );
  AOI22X1 U10963 ( .A0(n11667), .A1(n7937), .B0(n12883), .B1(n7887), .Y(n11666) );
  MX2X1 U10964 ( .A(n12881), .B(n11668), .S0(n11640), .Y(n11667) );
  AND2X1 U10965 ( .A(g25167), .B(n11669), .Y(n11640) );
  NAND2X1 U10966 ( .A(n12891), .B(n7458), .Y(n11668) );
  OAI21X1 U10967 ( .A0(n7938), .A1(n5351), .B0(n11670), .Y(n6049) );
  AOI22X1 U10968 ( .A0(n11159), .A1(n7733), .B0(n11160), .B1(n7304), .Y(n11670) );
  NAND2X1 U10969 ( .A(n11671), .B(n11672), .Y(n6048) );
  AOI22X1 U10970 ( .A0(n8456), .A1(n12891), .B0(n11673), .B1(n7938), .Y(n11672) );
  AOI22X1 U10971 ( .A0(n12877), .A1(n7910), .B0(n12881), .B1(test_se), .Y(
        n11671) );
  OAI21X1 U10972 ( .A0(n7865), .A1(n7691), .B0(n11674), .Y(n6047) );
  AOI22X1 U10973 ( .A0(n12880), .A1(n11675), .B0(n11643), .B1(n12879), .Y(
        n11674) );
  OAI21X1 U10974 ( .A0(test_se), .A1(n11676), .B0(n7920), .Y(n11675) );
  OAI21X1 U10975 ( .A0(n7921), .A1(n7232), .B0(n11677), .Y(n6046) );
  AOI21X1 U10976 ( .A0(n11643), .A1(n12878), .B0(n11678), .Y(n11677) );
  AOI21X1 U10977 ( .A0(n7865), .A1(n11634), .B0(n7511), .Y(n11678) );
  INVX1 U10978 ( .A(n11664), .Y(n11634) );
  NAND2X1 U10979 ( .A(n11679), .B(n11680), .Y(n6045) );
  MX2X1 U10980 ( .A(n7232), .B(n11654), .S0(n7853), .Y(n11680) );
  AOI22X1 U10981 ( .A0(n12890), .A1(n8456), .B0(n12891), .B1(n7873), .Y(n11679) );
  NOR2X1 U10982 ( .A(n8460), .B(n7972), .Y(n8456) );
  OAI22X1 U10983 ( .A0(n7865), .A1(n7529), .B0(n11681), .B1(n7972), .Y(n6044)
         );
  AOI22X1 U10984 ( .A0(n11682), .A1(n8460), .B0(n12889), .B1(n11683), .Y(
        n11681) );
  NOR2X1 U10985 ( .A(n12890), .B(n12891), .Y(n11682) );
  NAND2X1 U10986 ( .A(n11684), .B(n11685), .Y(n6043) );
  MX2X1 U10987 ( .A(n11686), .B(n11652), .S0(n11687), .Y(n11685) );
  NOR2X1 U10988 ( .A(n12889), .B(n11654), .Y(n11687) );
  NAND2X1 U10989 ( .A(n12891), .B(n8460), .Y(n11654) );
  NAND2X1 U10990 ( .A(n12884), .B(n7938), .Y(n11686) );
  AOI22X1 U10991 ( .A0(n7888), .A1(n7452), .B0(n12883), .B1(test_se), .Y(
        n11684) );
  NAND2X1 U10992 ( .A(n11688), .B(n11689), .Y(n6042) );
  AOI22X1 U10993 ( .A0(n11690), .A1(n12883), .B0(n11691), .B1(n11692), .Y(
        n11689) );
  INVX1 U10994 ( .A(n11683), .Y(n11692) );
  NAND2X1 U10995 ( .A(n12890), .B(n8460), .Y(n11683) );
  NOR2X1 U10996 ( .A(n7458), .B(n11652), .Y(n11691) );
  INVX1 U10997 ( .A(n11647), .Y(n11652) );
  AOI21X1 U10998 ( .A0(n7356), .A1(n11693), .B0(n7972), .Y(n11647) );
  AOI21X1 U10999 ( .A0(n11673), .A1(n12890), .B0(n7972), .Y(n11690) );
  AOI22X1 U11000 ( .A0(n12884), .A1(n7878), .B0(n12885), .B1(test_se), .Y(
        n11688) );
  NAND3X1 U11001 ( .A(n11694), .B(n11695), .C(n11696), .Y(n6041) );
  AOI22X1 U11002 ( .A0(n12887), .A1(n7909), .B0(n12889), .B1(test_se), .Y(
        n11696) );
  NAND3X1 U11003 ( .A(n11673), .B(g35), .C(n11697), .Y(n11695) );
  AOI21X1 U11004 ( .A0(n11693), .A1(n7356), .B0(n12891), .Y(n11697) );
  OAI21X1 U11005 ( .A0(n12891), .A1(n11698), .B0(n11642), .Y(n11694) );
  AND2X1 U11006 ( .A(n12888), .B(n7938), .Y(n11642) );
  INVX1 U11007 ( .A(n11673), .Y(n11698) );
  NOR2X1 U11008 ( .A(n7458), .B(n11659), .Y(n11673) );
  OAI21X1 U11009 ( .A0(n7865), .A1(n7590), .B0(n11699), .Y(n6040) );
  AOI21X1 U11010 ( .A0(n13015), .A1(n11700), .B0(n11701), .Y(n11699) );
  AOI21X1 U11011 ( .A0(n11702), .A1(n11703), .B0(n7314), .Y(n11701) );
  NAND3X1 U11012 ( .A(n11704), .B(n7617), .C(n7938), .Y(n11703) );
  OAI21X1 U11013 ( .A0(test_se), .A1(n11705), .B0(n7920), .Y(n11700) );
  AOI21X1 U11014 ( .A0(n11669), .A1(n7314), .B0(n11641), .Y(n11705) );
  INVX1 U11015 ( .A(n11706), .Y(n6039) );
  AOI22X1 U11016 ( .A0(n11707), .A1(n7938), .B0(n12874), .B1(n8593), .Y(n11706) );
  MX2X1 U11017 ( .A(n7602), .B(n11708), .S0(n11641), .Y(n11707) );
  NOR2X1 U11018 ( .A(n11704), .B(n11676), .Y(n11641) );
  NAND2X1 U11019 ( .A(n12879), .B(n7273), .Y(n11704) );
  XOR2X1 U11020 ( .A(n7314), .B(n7590), .Y(n11708) );
  OAI21X1 U11021 ( .A0(n12873), .A1(n7938), .B0(n11709), .Y(n6038) );
  MX2X1 U11022 ( .A(n11710), .B(n11711), .S0(n7591), .Y(n11709) );
  NAND2X1 U11023 ( .A(n11664), .B(n11635), .Y(n11711) );
  MX2X1 U11024 ( .A(n12871), .B(n12872), .S0(n11644), .Y(n6037) );
  OAI21X1 U11025 ( .A0(n11644), .A1(n7337), .B0(n11712), .Y(n6036) );
  MX2X1 U11026 ( .A(n11713), .B(n11714), .S0(n12871), .Y(n11712) );
  AOI21X1 U11027 ( .A0(n12872), .A1(n8461), .B0(n8593), .Y(n11714) );
  NAND3X1 U11028 ( .A(n7938), .B(n7591), .C(n8461), .Y(n11713) );
  OAI21X1 U11029 ( .A0(n11644), .A1(n7514), .B0(n11715), .Y(n6035) );
  MX2X1 U11030 ( .A(n11716), .B(n7337), .S0(n7958), .Y(n11715) );
  NAND2X1 U11031 ( .A(n8461), .B(n7514), .Y(n11716) );
  INVX1 U11032 ( .A(n11648), .Y(n11644) );
  NOR2X1 U11033 ( .A(n7972), .B(n8461), .Y(n11648) );
  NOR2X1 U11034 ( .A(n8462), .B(n11659), .Y(n8461) );
  INVX1 U11035 ( .A(n8460), .Y(n11659) );
  NAND3X1 U11036 ( .A(n11717), .B(n7356), .C(n8452), .Y(n8460) );
  INVX1 U11037 ( .A(g27831), .Y(n11717) );
  OR2X1 U11038 ( .A(n12889), .B(n12890), .Y(n8462) );
  OAI21X1 U11039 ( .A0(n8721), .A1(n7514), .B0(n11718), .Y(n6034) );
  AOI21X1 U11040 ( .A0(n12869), .A1(n11719), .B0(n11720), .Y(n11718) );
  INVX1 U11041 ( .A(n11710), .Y(n11719) );
  OAI21X1 U11042 ( .A0(n11710), .A1(n7239), .B0(n11721), .Y(n6033) );
  MX2X1 U11043 ( .A(n11722), .B(n11723), .S0(n12869), .Y(n11721) );
  NOR2X1 U11044 ( .A(n11720), .B(n8593), .Y(n11723) );
  INVX1 U11045 ( .A(n11724), .Y(n11720) );
  NAND3X1 U11046 ( .A(n11635), .B(n11669), .C(n12870), .Y(n11724) );
  NAND3X1 U11047 ( .A(n11635), .B(n7514), .C(n11664), .Y(n11722) );
  NOR2X1 U11048 ( .A(n11676), .B(n7972), .Y(n11664) );
  INVX1 U11049 ( .A(n11669), .Y(n11676) );
  NOR2X1 U11050 ( .A(n7273), .B(n7404), .Y(n11635) );
  AOI21X1 U11051 ( .A0(n7273), .A1(n7938), .B0(n11665), .Y(n11710) );
  OAI21X1 U11052 ( .A0(n12878), .A1(n7971), .B0(n11702), .Y(n11665) );
  INVX1 U11053 ( .A(n11643), .Y(n11702) );
  NOR2X1 U11054 ( .A(n7971), .B(n11669), .Y(n11643) );
  NOR2X1 U11055 ( .A(n11725), .B(n11554), .Y(n11669) );
  INVX1 U11056 ( .A(n11726), .Y(n11554) );
  AOI21X1 U11057 ( .A0(n13010), .A1(n11389), .B0(n11390), .Y(n11725) );
  OAI22X1 U11058 ( .A0(n7865), .A1(n7239), .B0(n11727), .B1(n7971), .Y(n6032)
         );
  AOI22X1 U11059 ( .A0(n11728), .A1(n11729), .B0(n12867), .B1(n11730), .Y(
        n11727) );
  NOR2X1 U11060 ( .A(n12866), .B(n12868), .Y(n11728) );
  MX2X1 U11061 ( .A(n12864), .B(n12853), .S0(n11731), .Y(n6031) );
  NAND2X1 U11062 ( .A(n11732), .B(n11733), .Y(n6030) );
  AOI22X1 U11063 ( .A0(n11734), .A1(n8450), .B0(n12865), .B1(n11735), .Y(
        n11733) );
  INVX1 U11064 ( .A(n11736), .Y(n11734) );
  AOI22X1 U11065 ( .A0(n12864), .A1(n7896), .B0(test_se), .B1(n7395), .Y(
        n11732) );
  NAND2X1 U11066 ( .A(n11737), .B(n11738), .Y(n6029) );
  MX2X1 U11067 ( .A(n11739), .B(n11736), .S0(n11740), .Y(n11738) );
  NOR2X1 U11068 ( .A(n12868), .B(n11741), .Y(n11740) );
  NAND2X1 U11069 ( .A(n12863), .B(n7938), .Y(n11739) );
  AOI22X1 U11070 ( .A0(n7907), .A1(n7395), .B0(n12865), .B1(test_se), .Y(
        n11737) );
  NAND2X1 U11071 ( .A(n11742), .B(n11743), .Y(n6028) );
  MX2X1 U11072 ( .A(n11744), .B(n11736), .S0(n11745), .Y(n11743) );
  NOR2X1 U11073 ( .A(n12866), .B(n11730), .Y(n11745) );
  NAND2X1 U11074 ( .A(n7938), .B(n7453), .Y(n11744) );
  AOI22X1 U11075 ( .A0(n12863), .A1(n7902), .B0(n12862), .B1(test_se), .Y(
        n11742) );
  NAND2X1 U11076 ( .A(n11746), .B(n11747), .Y(n6027) );
  AOI22X1 U11077 ( .A0(n11748), .A1(n11749), .B0(n12858), .B1(n11750), .Y(
        n11747) );
  NOR2X1 U11078 ( .A(n12856), .B(n11751), .Y(n11748) );
  AOI22X1 U11079 ( .A0(n12859), .A1(n7901), .B0(test_se), .B1(n7453), .Y(
        n11746) );
  OAI21X1 U11080 ( .A0(n7860), .A1(n7490), .B0(n11752), .Y(n6026) );
  AOI22X1 U11081 ( .A0(n11753), .A1(n7938), .B0(n12861), .B1(n7890), .Y(n11752) );
  MX2X1 U11082 ( .A(n11754), .B(n12859), .S0(n11755), .Y(n11753) );
  NAND2X1 U11083 ( .A(n12866), .B(n7405), .Y(n11754) );
  OAI21X1 U11084 ( .A0(n7860), .A1(n7686), .B0(n11756), .Y(n6025) );
  AOI22X1 U11085 ( .A0(n11757), .A1(n7938), .B0(n12855), .B1(n7892), .Y(n11756) );
  MX2X1 U11086 ( .A(n12866), .B(n12867), .S0(n11729), .Y(n11757) );
  NAND2X1 U11087 ( .A(n11758), .B(n11759), .Y(n6024) );
  MX2X1 U11088 ( .A(n11760), .B(n11761), .S0(n11762), .Y(n11759) );
  NOR2X1 U11089 ( .A(n7405), .B(n11763), .Y(n11762) );
  NAND2X1 U11090 ( .A(n11729), .B(n7470), .Y(n11763) );
  OAI21X1 U11091 ( .A0(n13038), .A1(n11589), .B0(g35), .Y(n11761) );
  NAND2X1 U11092 ( .A(n7938), .B(n7395), .Y(n11760) );
  AOI22X1 U11093 ( .A0(n12865), .A1(n7884), .B0(n12867), .B1(test_se), .Y(
        n11758) );
  OAI21X1 U11094 ( .A0(n7860), .A1(n7345), .B0(n11764), .Y(n6023) );
  AOI22X1 U11095 ( .A0(n12858), .A1(n11765), .B0(n11750), .B1(n12857), .Y(
        n11764) );
  OAI21X1 U11096 ( .A0(n11766), .A1(n11333), .B0(n7920), .Y(n11765) );
  INVX1 U11097 ( .A(n11365), .Y(n11333) );
  OAI21X1 U11098 ( .A0(n7921), .A1(n7208), .B0(n11767), .Y(n6022) );
  AOI21X1 U11099 ( .A0(n11750), .A1(n12856), .B0(n11768), .Y(n11767) );
  AOI21X1 U11100 ( .A0(n7860), .A1(n11769), .B0(n7555), .Y(n11768) );
  NAND2X1 U11101 ( .A(n11770), .B(n11771), .Y(n6021) );
  MX2X1 U11102 ( .A(n7208), .B(n11741), .S0(n7854), .Y(n11771) );
  AOI22X1 U11103 ( .A0(n11772), .A1(n8449), .B0(n12866), .B1(n7894), .Y(n11770) );
  AND2X1 U11104 ( .A(n7938), .B(n12868), .Y(n11772) );
  NAND2X1 U11105 ( .A(n11773), .B(n11774), .Y(n6020) );
  MX2X1 U11106 ( .A(n11775), .B(n11736), .S0(n11776), .Y(n11774) );
  NOR2X1 U11107 ( .A(n7405), .B(n11730), .Y(n11776) );
  NAND2X1 U11108 ( .A(n12868), .B(n11729), .Y(n11730) );
  NAND2X1 U11109 ( .A(n12861), .B(n7938), .Y(n11775) );
  AOI22X1 U11110 ( .A0(n12862), .A1(n7904), .B0(n12863), .B1(test_se), .Y(
        n11773) );
  NAND2X1 U11111 ( .A(n11777), .B(n11778), .Y(n6019) );
  MX2X1 U11112 ( .A(n11779), .B(n11736), .S0(n11780), .Y(n11778) );
  NOR2X1 U11113 ( .A(n12867), .B(n11741), .Y(n11780) );
  NAND2X1 U11114 ( .A(n12866), .B(n11729), .Y(n11741) );
  OAI21X1 U11115 ( .A0(n13038), .A1(n11589), .B0(n7922), .Y(n11736) );
  NAND2X1 U11116 ( .A(n8452), .B(g30332), .Y(n11589) );
  NAND2X1 U11117 ( .A(n12862), .B(n7938), .Y(n11779) );
  AOI22X1 U11118 ( .A0(n7895), .A1(n7453), .B0(n12861), .B1(test_se), .Y(
        n11777) );
  NAND3X1 U11119 ( .A(n11781), .B(n11782), .C(n11783), .Y(n6018) );
  AOI22X1 U11120 ( .A0(n12856), .A1(n7889), .B0(n12868), .B1(test_se), .Y(
        n11783) );
  NAND2X1 U11121 ( .A(n11750), .B(n13012), .Y(n11782) );
  AOI22X1 U11122 ( .A0(n11784), .A1(n11785), .B0(n11749), .B1(n11786), .Y(
        n11781) );
  NAND3X1 U11123 ( .A(n11787), .B(n11788), .C(n11789), .Y(n11786) );
  AOI22X1 U11124 ( .A0(n11751), .A1(n7395), .B0(n11790), .B1(n12865), .Y(
        n11789) );
  NAND3X1 U11125 ( .A(n7490), .B(n7292), .C(n12861), .Y(n11788) );
  OR2X1 U11126 ( .A(n12857), .B(n11791), .Y(n11787) );
  AOI22X1 U11127 ( .A0(n12863), .A1(n12856), .B0(n12858), .B1(n12862), .Y(
        n11791) );
  INVX1 U11128 ( .A(n11755), .Y(n11785) );
  NAND3X1 U11129 ( .A(n12857), .B(n7292), .C(n11792), .Y(n11755) );
  NOR2X1 U11130 ( .A(n12860), .B(n7971), .Y(n11784) );
  NAND2X1 U11131 ( .A(n11793), .B(n11794), .Y(n6017) );
  MX2X1 U11132 ( .A(n11795), .B(n11796), .S0(n7524), .Y(n11794) );
  NAND2X1 U11133 ( .A(n11797), .B(n7938), .Y(n11796) );
  AOI21X1 U11134 ( .A0(n11798), .A1(n11365), .B0(n7885), .Y(n11795) );
  NOR2X1 U11135 ( .A(n11388), .B(test_se), .Y(n11365) );
  NOR2X1 U11136 ( .A(n11766), .B(n11797), .Y(n11798) );
  NOR2X1 U11137 ( .A(n7522), .B(n11751), .Y(n11797) );
  AOI22X1 U11138 ( .A0(n12852), .A1(n11750), .B0(n12864), .B1(test_se), .Y(
        n11793) );
  OAI21X1 U11139 ( .A0(n8721), .A1(n7522), .B0(n11799), .Y(n6016) );
  AOI22X1 U11140 ( .A0(n11800), .A1(n11751), .B0(n11801), .B1(n7603), .Y(
        n11799) );
  OAI21X1 U11141 ( .A0(n11751), .A1(n7971), .B0(n11802), .Y(n11801) );
  INVX1 U11142 ( .A(n11750), .Y(n11802) );
  NOR2X1 U11143 ( .A(n7555), .B(n12858), .Y(n11751) );
  NOR2X1 U11144 ( .A(n11803), .B(n11769), .Y(n11800) );
  INVX1 U11145 ( .A(n11749), .Y(n11769) );
  XOR2X1 U11146 ( .A(n12864), .B(n7522), .Y(n11803) );
  OAI21X1 U11147 ( .A0(n12849), .A1(n7938), .B0(n11804), .Y(n6015) );
  MX2X1 U11148 ( .A(n11805), .B(n11806), .S0(n7592), .Y(n11804) );
  NAND2X1 U11149 ( .A(n11790), .B(n11749), .Y(n11806) );
  MX2X1 U11150 ( .A(n12847), .B(n12848), .S0(n11731), .Y(n6014) );
  OAI21X1 U11151 ( .A0(n11731), .A1(n7214), .B0(n11807), .Y(n6013) );
  MX2X1 U11152 ( .A(n11808), .B(n11809), .S0(n12847), .Y(n11807) );
  AOI21X1 U11153 ( .A0(n12848), .A1(n8450), .B0(n8593), .Y(n11809) );
  NAND3X1 U11154 ( .A(n7938), .B(n7592), .C(n8450), .Y(n11808) );
  OAI21X1 U11155 ( .A0(n11731), .A1(n7311), .B0(n11810), .Y(n6012) );
  MX2X1 U11156 ( .A(n11811), .B(n7214), .S0(n7959), .Y(n11810) );
  NAND2X1 U11157 ( .A(n8450), .B(n7311), .Y(n11811) );
  INVX1 U11158 ( .A(n11735), .Y(n11731) );
  NOR2X1 U11159 ( .A(n7971), .B(n8450), .Y(n11735) );
  NOR2X1 U11160 ( .A(n8448), .B(n8449), .Y(n8450) );
  INVX1 U11161 ( .A(n11729), .Y(n8449) );
  NAND3X1 U11162 ( .A(n11812), .B(n7367), .C(n8452), .Y(n11729) );
  INVX1 U11163 ( .A(n11813), .Y(n11812) );
  AOI21X1 U11164 ( .A0(n8244), .A1(n11814), .B0(n7912), .Y(n11813) );
  NOR2X1 U11165 ( .A(n7557), .B(n13053), .Y(n8244) );
  OR2X1 U11166 ( .A(n12867), .B(n12868), .Y(n8448) );
  OAI22X1 U11167 ( .A0(n11805), .A1(n7665), .B0(n11815), .B1(n7311), .Y(n6011)
         );
  AOI21X1 U11168 ( .A0(n11790), .A1(n11792), .B0(n8593), .Y(n11815) );
  OAI21X1 U11169 ( .A0(n11805), .A1(n7764), .B0(n11816), .Y(n6010) );
  MX2X1 U11170 ( .A(n11817), .B(n11818), .S0(n7665), .Y(n11816) );
  NAND3X1 U11171 ( .A(n11749), .B(n7311), .C(n11790), .Y(n11818) );
  NOR2X1 U11172 ( .A(n11819), .B(n7971), .Y(n11749) );
  AOI21X1 U11173 ( .A0(n11820), .A1(n12846), .B0(n8593), .Y(n11817) );
  NOR2X1 U11174 ( .A(n11819), .B(n11821), .Y(n11820) );
  INVX1 U11175 ( .A(n11792), .Y(n11819) );
  AOI21X1 U11176 ( .A0(n11821), .A1(n7938), .B0(n11750), .Y(n11805) );
  NOR2X1 U11177 ( .A(n7971), .B(n11792), .Y(n11750) );
  NOR2X1 U11178 ( .A(n11388), .B(n11766), .Y(n11792) );
  AOI21X1 U11179 ( .A0(n11389), .A1(n13008), .B0(n11390), .Y(n11766) );
  INVX1 U11180 ( .A(n11822), .Y(n11388) );
  INVX1 U11181 ( .A(n11790), .Y(n11821) );
  NOR2X1 U11182 ( .A(n7490), .B(n7292), .Y(n11790) );
  NAND3X1 U11183 ( .A(n11823), .B(n11824), .C(n11825), .Y(n6009) );
  NAND2X1 U11184 ( .A(n12845), .B(test_se), .Y(n11825) );
  NAND4X1 U11185 ( .A(n7938), .B(n11826), .C(n7510), .D(n7293), .Y(n11824) );
  NAND2X1 U11186 ( .A(n11827), .B(n11828), .Y(n11823) );
  MX2X1 U11187 ( .A(n12840), .B(n12826), .S0(n11829), .Y(n6008) );
  NAND2X1 U11188 ( .A(n11830), .B(n11831), .Y(n6007) );
  AOI22X1 U11189 ( .A0(n8435), .A1(n11832), .B0(n12841), .B1(n11833), .Y(
        n11831) );
  AOI22X1 U11190 ( .A0(n12840), .A1(n7874), .B0(test_se), .B1(n7396), .Y(
        n11830) );
  NAND2X1 U11191 ( .A(n11834), .B(n11835), .Y(n6006) );
  MX2X1 U11192 ( .A(n11836), .B(n11837), .S0(n11838), .Y(n11835) );
  NOR2X1 U11193 ( .A(n12844), .B(n11839), .Y(n11838) );
  NAND2X1 U11194 ( .A(n12839), .B(n7938), .Y(n11836) );
  AOI22X1 U11195 ( .A0(n7874), .A1(n7396), .B0(n12841), .B1(test_se), .Y(
        n11834) );
  NAND2X1 U11196 ( .A(n11840), .B(n11841), .Y(n6005) );
  MX2X1 U11197 ( .A(n11842), .B(n11837), .S0(n11843), .Y(n11841) );
  NOR2X1 U11198 ( .A(n12842), .B(n11828), .Y(n11843) );
  INVX1 U11199 ( .A(n11844), .Y(n11842) );
  AOI22X1 U11200 ( .A0(n12839), .A1(n7874), .B0(n12838), .B1(test_se), .Y(
        n11840) );
  NAND2X1 U11201 ( .A(n11845), .B(n11846), .Y(n6004) );
  AOI22X1 U11202 ( .A0(n11847), .A1(n11848), .B0(n12834), .B1(n11849), .Y(
        n11846) );
  NOR2X1 U11203 ( .A(n12832), .B(n11850), .Y(n11847) );
  AOI22X1 U11204 ( .A0(n12835), .A1(n7874), .B0(test_se), .B1(n7505), .Y(
        n11845) );
  OAI21X1 U11205 ( .A0(n7860), .A1(n7491), .B0(n11851), .Y(n6003) );
  AOI22X1 U11206 ( .A0(n11852), .A1(n7938), .B0(n12837), .B1(n7874), .Y(n11851) );
  MX2X1 U11207 ( .A(n11853), .B(n12835), .S0(n11854), .Y(n11852) );
  NAND2X1 U11208 ( .A(n12842), .B(n7257), .Y(n11853) );
  NAND2X1 U11209 ( .A(n11855), .B(n11856), .Y(n6002) );
  AOI22X1 U11210 ( .A0(n8431), .A1(n12842), .B0(n11827), .B1(n11826), .Y(
        n11856) );
  AOI22X1 U11211 ( .A0(n12831), .A1(n7874), .B0(n12835), .B1(test_se), .Y(
        n11855) );
  NAND2X1 U11212 ( .A(n11857), .B(n11858), .Y(n6001) );
  MX2X1 U11213 ( .A(n11859), .B(n11860), .S0(n11861), .Y(n11858) );
  NOR2X1 U11214 ( .A(n7257), .B(n11862), .Y(n11861) );
  NAND2X1 U11215 ( .A(n11826), .B(n7293), .Y(n11862) );
  OAI21X1 U11216 ( .A0(n13036), .A1(n11863), .B0(g35), .Y(n11860) );
  NAND2X1 U11217 ( .A(n7939), .B(n7396), .Y(n11859) );
  AOI22X1 U11218 ( .A0(n12841), .A1(n7874), .B0(n12843), .B1(test_se), .Y(
        n11857) );
  OAI21X1 U11219 ( .A0(n7860), .A1(n7692), .B0(n11864), .Y(n6000) );
  AOI22X1 U11220 ( .A0(n12834), .A1(n11865), .B0(n11849), .B1(n12833), .Y(
        n11864) );
  OAI21X1 U11221 ( .A0(n11866), .A1(n11433), .B0(n7920), .Y(n11865) );
  INVX1 U11222 ( .A(n11466), .Y(n11433) );
  OAI21X1 U11223 ( .A0(n7921), .A1(n7233), .B0(n11867), .Y(n5999) );
  AOI21X1 U11224 ( .A0(n11849), .A1(n12832), .B0(n11868), .Y(n11867) );
  AOI21X1 U11225 ( .A0(n7860), .A1(n11869), .B0(n7556), .Y(n11868) );
  NAND2X1 U11226 ( .A(n11870), .B(n11871), .Y(n5998) );
  MX2X1 U11227 ( .A(n7233), .B(n11839), .S0(n7853), .Y(n11871) );
  AOI22X1 U11228 ( .A0(n12844), .A1(n8431), .B0(n12842), .B1(n7874), .Y(n11870) );
  NOR2X1 U11229 ( .A(n11826), .B(n7971), .Y(n8431) );
  NAND2X1 U11230 ( .A(n11872), .B(n11873), .Y(n5997) );
  MX2X1 U11231 ( .A(n11874), .B(n11837), .S0(n11875), .Y(n11873) );
  NOR2X1 U11232 ( .A(n7257), .B(n11828), .Y(n11875) );
  NAND2X1 U11233 ( .A(n12844), .B(n11826), .Y(n11828) );
  INVX1 U11234 ( .A(n11832), .Y(n11837) );
  NAND2X1 U11235 ( .A(n12837), .B(n7939), .Y(n11874) );
  AOI22X1 U11236 ( .A0(n12838), .A1(n7874), .B0(n12839), .B1(test_se), .Y(
        n11872) );
  NAND3X1 U11237 ( .A(n11876), .B(n11877), .C(n11878), .Y(n5996) );
  AOI22X1 U11238 ( .A0(n7874), .A1(n7505), .B0(n12837), .B1(test_se), .Y(
        n11878) );
  NAND3X1 U11239 ( .A(n11832), .B(n7257), .C(n11879), .Y(n11877) );
  OAI21X1 U11240 ( .A0(n11693), .A1(n7971), .B0(n8438), .Y(n11832) );
  NAND2X1 U11241 ( .A(n13036), .B(n7939), .Y(n8438) );
  INVX1 U11242 ( .A(n11863), .Y(n11693) );
  NAND2X1 U11243 ( .A(n5529), .B(n8452), .Y(n11863) );
  NAND2X1 U11244 ( .A(n11880), .B(n12838), .Y(n11876) );
  INVX1 U11245 ( .A(n11881), .Y(n11880) );
  AOI21X1 U11246 ( .A0(n7939), .A1(n11839), .B0(n11827), .Y(n11881) );
  NOR2X1 U11247 ( .A(n7257), .B(n7971), .Y(n11827) );
  INVX1 U11248 ( .A(n11879), .Y(n11839) );
  NOR2X1 U11249 ( .A(n7293), .B(n8433), .Y(n11879) );
  OAI21X1 U11250 ( .A0(n7860), .A1(n7842), .B0(n11882), .Y(n5995) );
  AOI22X1 U11251 ( .A0(n7939), .A1(n11883), .B0(n12665), .B1(n7874), .Y(n11882) );
  NAND3X1 U11252 ( .A(n11884), .B(n11885), .C(n12666), .Y(n11883) );
  OAI21X1 U11253 ( .A0(n12666), .A1(n7860), .B0(n11886), .Y(n5994) );
  AOI21X1 U11254 ( .A0(n12664), .A1(n7874), .B0(n11887), .Y(n11886) );
  AOI21X1 U11255 ( .A0(n12663), .A1(n7758), .B0(n7971), .Y(n11887) );
  OAI21X1 U11256 ( .A0(n7860), .A1(n7352), .B0(n11888), .Y(n5993) );
  AOI22X1 U11257 ( .A0(n12661), .A1(n8108), .B0(g37), .B1(n7939), .Y(n11888)
         );
  MX2X1 U11258 ( .A(g37), .B(n7684), .S0(n7853), .Y(n5992) );
  OAI21X1 U11259 ( .A0(n7860), .A1(n7597), .B0(n11889), .Y(n5991) );
  AOI22X1 U11260 ( .A0(n11890), .A1(n12453), .B0(n7874), .B1(g18881), .Y(
        n11889) );
  NOR2X1 U11261 ( .A(n12450), .B(n8140), .Y(n11890) );
  NAND4X1 U11262 ( .A(n12541), .B(n7939), .C(n12540), .D(n11891), .Y(n8140) );
  NOR2X1 U11263 ( .A(n7353), .B(n11892), .Y(n11891) );
  NAND2X1 U11264 ( .A(n12452), .B(n12539), .Y(n11892) );
  OAI21X1 U11265 ( .A0(n7860), .A1(n7822), .B0(n11893), .Y(n5990) );
  AOI21X1 U11266 ( .A0(n12410), .A1(n11894), .B0(n8163), .Y(n11893) );
  NOR2X1 U11267 ( .A(n7759), .B(n7971), .Y(n8163) );
  NAND2X1 U11268 ( .A(n7921), .B(n11895), .Y(n11894) );
  NAND4X1 U11269 ( .A(n12411), .B(n12413), .C(n12412), .D(n7860), .Y(n11895)
         );
  MX2X1 U11270 ( .A(n12676), .B(g10306), .S0(n7852), .Y(n5989) );
  OAI21X1 U11271 ( .A0(n7860), .A1(n7734), .B0(n11896), .Y(n5988) );
  AOI22X1 U11272 ( .A0(n12433), .A1(n11897), .B0(n7939), .B1(n11898), .Y(
        n11896) );
  OAI21X1 U11273 ( .A0(n12433), .A1(n7616), .B0(n11899), .Y(n11898) );
  XOR2X1 U11274 ( .A(n12436), .B(n7632), .Y(n11899) );
  OAI21X1 U11275 ( .A0(test_se), .A1(n12438), .B0(n7920), .Y(n11897) );
  INVX1 U11276 ( .A(n11900), .Y(n5987) );
  AOI21X1 U11277 ( .A0(n12429), .A1(n7860), .B0(n11901), .Y(n11900) );
  AOI21X1 U11278 ( .A0(n7860), .A1(n11902), .B0(n7815), .Y(n11901) );
  NAND3X1 U11279 ( .A(g35), .B(n7263), .C(n11903), .Y(n11902) );
  INVX1 U11280 ( .A(n11904), .Y(n11903) );
  INVX1 U11281 ( .A(n11905), .Y(n5986) );
  AOI22X1 U11282 ( .A0(n12441), .A1(n7939), .B0(n12432), .B1(test_se), .Y(
        n11905) );
  OAI21X1 U11283 ( .A0(n5305), .A1(n7860), .B0(n11906), .Y(n5985) );
  AOI22X1 U11284 ( .A0(n8168), .A1(n8196), .B0(n12430), .B1(n8170), .Y(n11906)
         );
  OAI21X1 U11285 ( .A0(test_se), .A1(n7475), .B0(n7920), .Y(n8170) );
  NOR2X1 U11286 ( .A(n7970), .B(n7263), .Y(n8168) );
  INVX1 U11287 ( .A(n11907), .Y(n5984) );
  MX2X1 U11288 ( .A(n7683), .B(n5304), .S0(n7853), .Y(n11907) );
  INVX1 U11289 ( .A(n11908), .Y(n5983) );
  MX2X1 U11290 ( .A(n5304), .B(n5305), .S0(n7852), .Y(n11908) );
  OAI21X1 U11291 ( .A0(n7860), .A1(n7843), .B0(n11909), .Y(n5982) );
  OAI21X1 U11292 ( .A0(n12428), .A1(n7530), .B0(n7922), .Y(n11909) );
  OAI22X1 U11293 ( .A0(n7860), .A1(n7633), .B0(n11910), .B1(n7317), .Y(n5981)
         );
  AOI21X1 U11294 ( .A0(n11911), .A1(n7860), .B0(n7879), .Y(n11910) );
  NAND3X1 U11295 ( .A(n7228), .B(n7530), .C(n7245), .Y(n11911) );
  NAND3X1 U11296 ( .A(n11912), .B(n7921), .C(n12428), .Y(n5980) );
  NAND3X1 U11297 ( .A(n12449), .B(n7860), .C(n12427), .Y(n11912) );
  OAI21X1 U11298 ( .A0(n7860), .A1(n7530), .B0(n11913), .Y(n5979) );
  AOI22X1 U11299 ( .A0(n7939), .A1(n11914), .B0(n12537), .B1(n7914), .Y(n11913) );
  OAI21X1 U11300 ( .A0(n7317), .A1(n7228), .B0(n7633), .Y(n11914) );
  OAI21X1 U11301 ( .A0(n7860), .A1(n7762), .B0(n11915), .Y(n5978) );
  AOI22X1 U11302 ( .A0(n12448), .A1(n7886), .B0(n12449), .B1(n7939), .Y(n11915) );
  OAI21X1 U11303 ( .A0(n7939), .A1(n5297), .B0(n11916), .Y(n5977) );
  OR2X1 U11304 ( .A(n11917), .B(n8158), .Y(n5976) );
  MX2X1 U11305 ( .A(n12424), .B(n12423), .S0(n7853), .Y(n11917) );
  NAND2X1 U11306 ( .A(n5293), .B(n8155), .Y(n5975) );
  NAND2X1 U11307 ( .A(n5292), .B(n8155), .Y(n5974) );
  NAND2X1 U11308 ( .A(n11918), .B(n11919), .Y(n5973) );
  MX2X1 U11309 ( .A(n11920), .B(n11921), .S0(n7597), .Y(n11919) );
  NAND2X1 U11310 ( .A(n11922), .B(n8162), .Y(n11921) );
  AOI21X1 U11311 ( .A0(n11922), .A1(n11923), .B0(n7875), .Y(n11920) );
  AOI22X1 U11312 ( .A0(n11924), .A1(n12447), .B0(n12417), .B1(test_se), .Y(
        n11918) );
  NOR2X1 U11313 ( .A(n12418), .B(n7970), .Y(n11924) );
  OAI21X1 U11314 ( .A0(n7860), .A1(n7844), .B0(n11925), .Y(n5972) );
  AOI22X1 U11315 ( .A0(n12675), .A1(n7876), .B0(n12441), .B1(n7939), .Y(n11925) );
  NAND2X1 U11316 ( .A(n11926), .B(n11927), .Y(n5971) );
  AOI21X1 U11317 ( .A0(n7939), .A1(n11928), .B0(n11929), .Y(n11927) );
  NAND2X1 U11318 ( .A(n11930), .B(n11931), .Y(n11928) );
  NAND3X1 U11319 ( .A(n12815), .B(n11932), .C(n12437), .Y(n11931) );
  AOI22X1 U11320 ( .A0(n12438), .A1(n7908), .B0(test_se), .B1(n7275), .Y(
        n11926) );
  OAI21X1 U11321 ( .A0(n7859), .A1(n7475), .B0(n11933), .Y(n5970) );
  AOI21X1 U11322 ( .A0(n12817), .A1(n7939), .B0(n11934), .Y(n11933) );
  AOI21X1 U11323 ( .A0(n7921), .A1(n11935), .B0(n7738), .Y(n11934) );
  NAND3X1 U11324 ( .A(n12814), .B(n7859), .C(n8169), .Y(n11935) );
  NAND2X1 U11325 ( .A(n11936), .B(n11937), .Y(n5969) );
  NAND3X1 U11326 ( .A(n12438), .B(n8169), .C(n11938), .Y(n11937) );
  MX2X1 U11327 ( .A(n7263), .B(n7760), .S0(n7853), .Y(n11936) );
  MX2X1 U11328 ( .A(n12436), .B(g7243), .S0(n7853), .Y(n5968) );
  NAND2X1 U11329 ( .A(n11939), .B(n11940), .Y(n5967) );
  AOI21X1 U11330 ( .A0(n11938), .A1(n8169), .B0(n11929), .Y(n11940) );
  INVX1 U11331 ( .A(n11941), .Y(n11929) );
  NAND3X1 U11332 ( .A(n7275), .B(n7475), .C(n7939), .Y(n11941) );
  AOI22X1 U11333 ( .A0(n12817), .A1(n7915), .B0(n12816), .B1(test_se), .Y(
        n11939) );
  MX2X1 U11334 ( .A(g7243), .B(g7257), .S0(n7852), .Y(n5966) );
  INVX1 U11335 ( .A(n11942), .Y(n5965) );
  AOI22X1 U11336 ( .A0(n12437), .A1(n7882), .B0(test_se), .B1(g7257), .Y(
        n11942) );
  OAI21X1 U11337 ( .A0(n7859), .A1(n7616), .B0(n11943), .Y(n5964) );
  AOI22X1 U11338 ( .A0(n7939), .A1(n8166), .B0(n12813), .B1(n8108), .Y(n11943)
         );
  OAI21X1 U11339 ( .A0(n8169), .A1(n7263), .B0(n11930), .Y(n8166) );
  NAND3X1 U11340 ( .A(n7263), .B(n7761), .C(n8169), .Y(n11930) );
  NOR2X1 U11341 ( .A(n7275), .B(n11932), .Y(n8169) );
  NAND4X1 U11342 ( .A(n5289), .B(n5285), .C(n7344), .D(n7760), .Y(n11932) );
  INVX1 U11343 ( .A(n11944), .Y(n5963) );
  AOI21X1 U11344 ( .A0(n8196), .A1(n11938), .B0(n11945), .Y(n11944) );
  INVX1 U11345 ( .A(n11946), .Y(n11945) );
  MX2X1 U11346 ( .A(n11947), .B(n12431), .S0(n7958), .Y(n11946) );
  NAND2X1 U11347 ( .A(n12430), .B(n7475), .Y(n11947) );
  NOR2X1 U11348 ( .A(n7970), .B(n12814), .Y(n11938) );
  NOR2X1 U11349 ( .A(n11904), .B(n12429), .Y(n8196) );
  NAND4X1 U11350 ( .A(n12431), .B(n5305), .C(n5304), .D(n7683), .Y(n11904) );
  MX2X1 U11351 ( .A(g12832), .B(n7684), .S0(n7853), .Y(n5962) );
  OAI21X1 U11352 ( .A0(n7859), .A1(n7761), .B0(n11948), .Y(n5961) );
  MX2X1 U11353 ( .A(n11949), .B(n11950), .S0(n12434), .Y(n11948) );
  AOI21X1 U11354 ( .A0(n5311), .A1(n7859), .B0(n7891), .Y(n11950) );
  NAND2X1 U11355 ( .A(n7939), .B(g10306), .Y(n11949) );
  NAND2X1 U11356 ( .A(n11951), .B(n11952), .Y(n5960) );
  AOI21X1 U11357 ( .A0(n12417), .A1(n7873), .B0(n8157), .Y(n11952) );
  AOI22X1 U11358 ( .A0(n7939), .A1(n7822), .B0(n12416), .B1(test_se), .Y(
        n11951) );
  OAI21X1 U11359 ( .A0(n8150), .A1(n11953), .B0(n11954), .Y(n5959) );
  OAI21X1 U11360 ( .A0(n8593), .A1(n11955), .B0(n7456), .Y(n11954) );
  XOR2X1 U11361 ( .A(n12422), .B(n8162), .Y(n11955) );
  INVX1 U11362 ( .A(n11923), .Y(n8162) );
  NAND4X1 U11363 ( .A(n12419), .B(n12420), .C(n12421), .D(n12424), .Y(n11923)
         );
  INVX1 U11364 ( .A(n11922), .Y(n11953) );
  NOR2X1 U11365 ( .A(n7456), .B(n7970), .Y(n11922) );
  INVX1 U11366 ( .A(n8588), .Y(n8150) );
  NAND2X1 U11367 ( .A(n11956), .B(n11957), .Y(n8588) );
  NAND3X1 U11368 ( .A(n11958), .B(n12444), .C(n11959), .Y(n11957) );
  XOR2X1 U11369 ( .A(n7359), .B(n12445), .Y(n11959) );
  XOR2X1 U11370 ( .A(n12443), .B(n7355), .Y(n11958) );
  MX2X1 U11371 ( .A(n11960), .B(n11961), .S0(n7355), .Y(n11956) );
  NAND3X1 U11372 ( .A(n12445), .B(n7359), .C(n12443), .Y(n11961) );
  OR2X1 U11373 ( .A(n7359), .B(n12445), .Y(n11960) );
  NAND2X1 U11374 ( .A(n11962), .B(n11916), .Y(n5958) );
  AOI21X1 U11375 ( .A0(n8157), .A1(n12440), .B0(n8158), .Y(n11916) );
  NOR2X1 U11376 ( .A(n7970), .B(n12425), .Y(n8157) );
  AOI22X1 U11377 ( .A0(n12441), .A1(n7873), .B0(test_se), .B1(g10306), .Y(
        n11962) );
  NAND2X1 U11378 ( .A(n5281), .B(n8155), .Y(n5957) );
  INVX1 U11379 ( .A(n8158), .Y(n8155) );
  OR2X1 U11380 ( .A(n11963), .B(n8158), .Y(n5956) );
  MX2X1 U11381 ( .A(n12409), .B(n12408), .S0(n7852), .Y(n11963) );
  MX2X1 U11382 ( .A(g18096), .B(n12411), .S0(n7959), .Y(n5955) );
  OR2X1 U11383 ( .A(n11964), .B(n8158), .Y(n5954) );
  NOR2X1 U11384 ( .A(n7685), .B(n7970), .Y(n8158) );
  MX2X1 U11385 ( .A(n12410), .B(n12409), .S0(n7852), .Y(n11964) );
  NAND3X1 U11386 ( .A(n11965), .B(n11966), .C(n11967), .Y(n5953) );
  AOI22X1 U11387 ( .A0(n12832), .A1(n7873), .B0(n12844), .B1(test_se), .Y(
        n11967) );
  NAND2X1 U11388 ( .A(n11849), .B(n13014), .Y(n11966) );
  AOI22X1 U11389 ( .A0(n11968), .A1(n11844), .B0(n11848), .B1(n11969), .Y(
        n11965) );
  NAND3X1 U11390 ( .A(n11970), .B(n11971), .C(n11972), .Y(n11969) );
  AOI22X1 U11391 ( .A0(n11850), .A1(n7396), .B0(n11973), .B1(n12841), .Y(
        n11972) );
  NAND3X1 U11392 ( .A(n7491), .B(n7294), .C(n12837), .Y(n11971) );
  OR2X1 U11393 ( .A(n12833), .B(n11974), .Y(n11970) );
  AOI22X1 U11394 ( .A0(n12839), .A1(n12832), .B0(n12834), .B1(n12838), .Y(
        n11974) );
  NOR2X1 U11395 ( .A(n7970), .B(n12836), .Y(n11844) );
  INVX1 U11396 ( .A(n11854), .Y(n11968) );
  NAND3X1 U11397 ( .A(n12833), .B(n7294), .C(n11975), .Y(n11854) );
  NAND2X1 U11398 ( .A(n11976), .B(n11977), .Y(n5952) );
  MX2X1 U11399 ( .A(n11978), .B(n11979), .S0(n7324), .Y(n11977) );
  NAND2X1 U11400 ( .A(n11980), .B(n7939), .Y(n11979) );
  AOI21X1 U11401 ( .A0(n11981), .A1(n11466), .B0(n7873), .Y(n11978) );
  NOR2X1 U11402 ( .A(n11489), .B(test_se), .Y(n11466) );
  NOR2X1 U11403 ( .A(n11866), .B(n11980), .Y(n11981) );
  NOR2X1 U11404 ( .A(n7523), .B(n11850), .Y(n11980) );
  AOI22X1 U11405 ( .A0(n12825), .A1(n11849), .B0(n12840), .B1(test_se), .Y(
        n11976) );
  OAI21X1 U11406 ( .A0(n8721), .A1(n7523), .B0(n11982), .Y(n5951) );
  AOI22X1 U11407 ( .A0(n11983), .A1(n11850), .B0(n11984), .B1(n7604), .Y(
        n11982) );
  OAI21X1 U11408 ( .A0(n11850), .A1(n7970), .B0(n11985), .Y(n11984) );
  INVX1 U11409 ( .A(n11849), .Y(n11985) );
  NOR2X1 U11410 ( .A(n7556), .B(n12834), .Y(n11850) );
  NOR2X1 U11411 ( .A(n11986), .B(n11869), .Y(n11983) );
  INVX1 U11412 ( .A(n11848), .Y(n11869) );
  XOR2X1 U11413 ( .A(n12840), .B(n7523), .Y(n11986) );
  OAI21X1 U11414 ( .A0(n12824), .A1(n7939), .B0(n11987), .Y(n5950) );
  MX2X1 U11415 ( .A(n11988), .B(n11989), .S0(n7593), .Y(n11987) );
  NAND2X1 U11416 ( .A(n11973), .B(n11848), .Y(n11989) );
  MX2X1 U11417 ( .A(n12822), .B(n12823), .S0(n11829), .Y(n5949) );
  OAI21X1 U11418 ( .A0(n11829), .A1(n7649), .B0(n11990), .Y(n5948) );
  MX2X1 U11419 ( .A(n11991), .B(n11992), .S0(n12822), .Y(n11990) );
  AOI21X1 U11420 ( .A0(n12823), .A1(n8435), .B0(n8593), .Y(n11992) );
  NAND3X1 U11421 ( .A(n7939), .B(n7593), .C(n8435), .Y(n11991) );
  OAI21X1 U11422 ( .A0(n11829), .A1(n7312), .B0(n11993), .Y(n5947) );
  MX2X1 U11423 ( .A(n11994), .B(n7649), .S0(n7960), .Y(n11993) );
  NAND2X1 U11424 ( .A(n8435), .B(n7312), .Y(n11994) );
  INVX1 U11425 ( .A(n11833), .Y(n11829) );
  NOR2X1 U11426 ( .A(n7970), .B(n8435), .Y(n11833) );
  NOR2X1 U11427 ( .A(n8439), .B(n8433), .Y(n8435) );
  INVX1 U11428 ( .A(n11826), .Y(n8433) );
  NAND3X1 U11429 ( .A(n11995), .B(n7282), .C(n8452), .Y(n11826) );
  AND2X1 U11430 ( .A(n8779), .B(n8784), .Y(n8452) );
  NOR2X1 U11431 ( .A(n7244), .B(n12892), .Y(n8779) );
  INVX1 U11432 ( .A(n11996), .Y(n11995) );
  AOI21X1 U11433 ( .A0(n11814), .A1(n8691), .B0(n7933), .Y(n11996) );
  INVX1 U11434 ( .A(n8690), .Y(n8691) );
  NAND2X1 U11435 ( .A(n13053), .B(n13054), .Y(n8690) );
  NAND2X1 U11436 ( .A(n7257), .B(n7510), .Y(n8439) );
  OAI22X1 U11437 ( .A0(n11988), .A1(n7666), .B0(n11997), .B1(n7312), .Y(n5946)
         );
  AOI21X1 U11438 ( .A0(n11973), .A1(n11975), .B0(n8593), .Y(n11997) );
  OAI21X1 U11439 ( .A0(n11988), .A1(n7338), .B0(n11998), .Y(n5945) );
  MX2X1 U11440 ( .A(n11999), .B(n12000), .S0(n7666), .Y(n11998) );
  NAND3X1 U11441 ( .A(n11848), .B(n7312), .C(n11973), .Y(n12000) );
  NOR2X1 U11442 ( .A(n12001), .B(n7970), .Y(n11848) );
  AOI21X1 U11443 ( .A0(n12002), .A1(n12821), .B0(n8593), .Y(n11999) );
  INVX1 U11444 ( .A(n8721), .Y(n8593) );
  NOR2X1 U11445 ( .A(n12001), .B(n12003), .Y(n12002) );
  INVX1 U11446 ( .A(n11975), .Y(n12001) );
  AOI21X1 U11447 ( .A0(n12003), .A1(n7939), .B0(n11849), .Y(n11988) );
  NOR2X1 U11448 ( .A(n7970), .B(n11975), .Y(n11849) );
  NOR2X1 U11449 ( .A(n11489), .B(n11866), .Y(n11975) );
  AOI21X1 U11450 ( .A0(n11389), .A1(n13011), .B0(n11390), .Y(n11866) );
  INVX1 U11451 ( .A(n12004), .Y(n11390) );
  INVX1 U11452 ( .A(n12005), .Y(n11389) );
  NAND3X1 U11453 ( .A(n12006), .B(n7319), .C(n13026), .Y(n12005) );
  INVX1 U11454 ( .A(n12007), .Y(n11489) );
  INVX1 U11455 ( .A(n11973), .Y(n12003) );
  NOR2X1 U11456 ( .A(n7491), .B(n7294), .Y(n11973) );
  NAND2X1 U11457 ( .A(n12008), .B(n12009), .Y(n5944) );
  AOI22X1 U11458 ( .A0(n11159), .A1(n7686), .B0(n11160), .B1(n7303), .Y(n12009) );
  AOI22X1 U11459 ( .A0(n7873), .A1(n7304), .B0(test_se), .B1(n7377), .Y(n12008) );
  OAI21X1 U11460 ( .A0(n12699), .A1(n7939), .B0(n12010), .Y(n5943) );
  AOI22X1 U11461 ( .A0(n11159), .A1(n7687), .B0(n12698), .B1(n11160), .Y(
        n12010) );
  NAND2X1 U11462 ( .A(n12011), .B(n12012), .Y(n5942) );
  AOI22X1 U11463 ( .A0(n11159), .A1(n7735), .B0(n11160), .B1(n7329), .Y(n12012) );
  AOI22X1 U11464 ( .A0(n7873), .A1(n7305), .B0(test_se), .B1(n7218), .Y(n12011) );
  OAI21X1 U11465 ( .A0(n12687), .A1(n7940), .B0(n12013), .Y(n5941) );
  AOI22X1 U11466 ( .A0(n11159), .A1(n7736), .B0(n11160), .B1(n7306), .Y(n12013) );
  INVX1 U11467 ( .A(n12014), .Y(n11159) );
  NAND3X1 U11468 ( .A(n11626), .B(n12015), .C(n11160), .Y(n12014) );
  AOI21X1 U11469 ( .A0(n12006), .A1(n13031), .B0(n7970), .Y(n11160) );
  INVX1 U11470 ( .A(n12006), .Y(n12015) );
  NAND4X1 U11471 ( .A(n13029), .B(n13030), .C(n13031), .D(n13026), .Y(n11626)
         );
  OAI21X1 U11472 ( .A0(n12686), .A1(n7859), .B0(n12016), .Y(n5940) );
  AOI22X1 U11473 ( .A0(n7940), .A1(n8179), .B0(n7873), .B1(n7297), .Y(n12016)
         );
  INVX1 U11474 ( .A(n12017), .Y(n8179) );
  MX2X1 U11475 ( .A(n12018), .B(n12019), .S0(n12020), .Y(n12017) );
  NAND2X1 U11476 ( .A(n12021), .B(n12022), .Y(n12019) );
  AOI22X1 U11477 ( .A0(n11822), .A1(n7524), .B0(n11618), .B1(n7315), .Y(n12022) );
  AOI22X1 U11478 ( .A0(n12007), .A1(n7324), .B0(n11726), .B1(n7617), .Y(n12021) );
  NAND2X1 U11479 ( .A(n12023), .B(n12024), .Y(n12018) );
  AOI22X1 U11480 ( .A0(n11822), .A1(n7377), .B0(n13009), .B1(n11618), .Y(
        n12024) );
  AOI22X1 U11481 ( .A0(n12007), .A1(n7414), .B0(n11726), .B1(n7297), .Y(n12023) );
  OAI21X1 U11482 ( .A0(n7859), .A1(g30331), .B0(n12025), .Y(n5939) );
  AOI22X1 U11483 ( .A0(n7940), .A1(n8181), .B0(n7873), .B1(n7381), .Y(n12025)
         );
  INVX1 U11484 ( .A(n12026), .Y(n8181) );
  MX2X1 U11485 ( .A(n12027), .B(n12028), .S0(n12020), .Y(n12026) );
  NAND4X1 U11486 ( .A(n12004), .B(n12006), .C(n7319), .D(n7688), .Y(n12020) );
  NOR2X1 U11487 ( .A(n13029), .B(n13030), .Y(n12006) );
  NAND2X1 U11488 ( .A(n12029), .B(n12030), .Y(n12028) );
  AOI22X1 U11489 ( .A0(n11822), .A1(n7594), .B0(n11618), .B1(n7325), .Y(n12030) );
  AOI22X1 U11490 ( .A0(n12007), .A1(n7595), .B0(n11726), .B1(n7326), .Y(n12029) );
  NAND2X1 U11491 ( .A(n12031), .B(n12032), .Y(n12027) );
  AOI22X1 U11492 ( .A0(n11822), .A1(n7378), .B0(n11618), .B1(n7218), .Y(n12032) );
  NOR2X1 U11493 ( .A(n7574), .B(n7320), .Y(n11618) );
  NOR2X1 U11494 ( .A(n7320), .B(n13033), .Y(n11822) );
  AOI22X1 U11495 ( .A0(n12007), .A1(n7271), .B0(n11726), .B1(n7381), .Y(n12031) );
  NOR2X1 U11496 ( .A(n13032), .B(n13033), .Y(n11726) );
  NOR2X1 U11497 ( .A(n7574), .B(n13032), .Y(n12007) );
  INVX1 U11498 ( .A(n12033), .Y(n5938) );
  AOI22X1 U11499 ( .A0(n8562), .A1(n12034), .B0(n12241), .B1(n7970), .Y(n12033) );
  XOR2X1 U11500 ( .A(n12227), .B(n12035), .Y(n12034) );
  OAI21X1 U11501 ( .A0(n7940), .A1(n7695), .B0(n12036), .Y(n5937) );
  MX2X1 U11502 ( .A(n12037), .B(n12226), .S0(n12038), .Y(n12036) );
  NAND2X1 U11503 ( .A(n8562), .B(n12226), .Y(n12037) );
  OAI21X1 U11504 ( .A0(n8721), .A1(n7737), .B0(n12039), .Y(n5936) );
  MX2X1 U11505 ( .A(n12040), .B(n12225), .S0(n10945), .Y(n12039) );
  AND2X1 U11506 ( .A(n12226), .B(n12038), .Y(n10945) );
  NOR2X1 U11507 ( .A(n12041), .B(n7695), .Y(n12038) );
  OAI21X1 U11508 ( .A0(n671), .A1(n12241), .B0(n12035), .Y(n12041) );
  AOI21X1 U11509 ( .A0(g12184), .A1(n671), .B0(n10980), .Y(n12035) );
  NAND2X1 U11510 ( .A(n12042), .B(n12043), .Y(n10980) );
  MX2X1 U11511 ( .A(n12044), .B(n12045), .S0(n7385), .Y(n12043) );
  NAND2X1 U11512 ( .A(n12921), .B(n7251), .Y(n12045) );
  NAND2X1 U11513 ( .A(n12923), .B(n7463), .Y(n12044) );
  AOI21X1 U11514 ( .A0(n12924), .A1(n12925), .B0(n10914), .Y(n12042) );
  NAND2X1 U11515 ( .A(n8562), .B(n12225), .Y(n12040) );
  INVX1 U11516 ( .A(n10948), .Y(n8562) );
  OAI21X1 U11517 ( .A0(n12241), .A1(n671), .B0(n7922), .Y(n10948) );
  NOR2X1 U11518 ( .A(test_se), .B(n7873), .Y(n8721) );
  OAI21X1 U11519 ( .A0(n7859), .A1(n7639), .B0(n12046), .Y(n5935) );
  AOI22X1 U11520 ( .A0(n12047), .A1(n7940), .B0(n12159), .B1(n12048), .Y(
        n12046) );
  OAI21X1 U11521 ( .A0(test_se), .A1(n10914), .B0(n7920), .Y(n12048) );
  AND2X1 U11522 ( .A(n7385), .B(n10914), .Y(n12047) );
  NAND3X1 U11523 ( .A(n12049), .B(n12050), .C(n11084), .Y(n10914) );
  INVX1 U11524 ( .A(n11019), .Y(n11084) );
  OAI21X1 U11525 ( .A0(n7859), .A1(n7816), .B0(n12051), .Y(n5934) );
  AOI22X1 U11526 ( .A0(n10853), .A1(n12850), .B0(n12186), .B1(n8211), .Y(
        n12051) );
  NAND2X1 U11527 ( .A(n12052), .B(n12053), .Y(n5933) );
  AOI22X1 U11528 ( .A0(n10853), .A1(n12178), .B0(n12177), .B1(n8211), .Y(
        n12053) );
  NOR2X1 U11529 ( .A(n12054), .B(n7969), .Y(n10853) );
  AOI22X1 U11530 ( .A0(n7873), .A1(n7454), .B0(n12186), .B1(test_se), .Y(
        n12052) );
  MX2X1 U11531 ( .A(n12177), .B(n12921), .S0(n8211), .Y(n5932) );
  OAI21X1 U11532 ( .A0(n7859), .A1(n7463), .B0(n12055), .Y(n5931) );
  AOI22X1 U11533 ( .A0(n8210), .A1(n7251), .B0(n8211), .B1(n12171), .Y(n12055)
         );
  NAND2X1 U11534 ( .A(n12056), .B(n12057), .Y(n5930) );
  MX2X1 U11535 ( .A(n12058), .B(n12059), .S0(n7540), .Y(n12057) );
  NAND2X1 U11536 ( .A(n12060), .B(n10848), .Y(n12059) );
  NAND2X1 U11537 ( .A(n10841), .B(n12061), .Y(n12058) );
  INVX1 U11538 ( .A(n12060), .Y(n12061) );
  NOR2X1 U11539 ( .A(n10849), .B(n7525), .Y(n12060) );
  INVX1 U11540 ( .A(n10847), .Y(n10849) );
  NOR2X1 U11541 ( .A(n7696), .B(n8116), .Y(n10847) );
  AND2X1 U11542 ( .A(n10848), .B(n7940), .Y(n10841) );
  AOI21X1 U11543 ( .A0(n10843), .A1(n10837), .B0(n7407), .Y(n10848) );
  INVX1 U11544 ( .A(n12062), .Y(n10837) );
  NAND4X1 U11545 ( .A(n12178), .B(n12063), .C(n12064), .D(n12065), .Y(n12062)
         );
  NOR2X1 U11546 ( .A(n12186), .B(n12066), .Y(n12065) );
  OR2X1 U11547 ( .A(n12179), .B(n12177), .Y(n12066) );
  XOR2X1 U11548 ( .A(n7535), .B(n12169), .Y(n12064) );
  XOR2X1 U11549 ( .A(n7463), .B(n7251), .Y(n12063) );
  INVX1 U11550 ( .A(n8116), .Y(n10843) );
  NAND4X1 U11551 ( .A(n12067), .B(n12926), .C(n12068), .D(n7284), .Y(n8116) );
  NOR2X1 U11552 ( .A(n12267), .B(n12928), .Y(n12068) );
  NOR2X1 U11553 ( .A(n10870), .B(n7462), .Y(n12067) );
  NAND3X1 U11554 ( .A(n12069), .B(n12932), .C(n12931), .Y(n10870) );
  AOI22X1 U11555 ( .A0(n12168), .A1(n7873), .B0(n12490), .B1(test_se), .Y(
        n12056) );
  OAI21X1 U11556 ( .A0(n7867), .A1(n7540), .B0(n12070), .Y(n5929) );
  AOI22X1 U11557 ( .A0(n12921), .A1(n8210), .B0(n8211), .B1(n7251), .Y(n12070)
         );
  NOR2X1 U11558 ( .A(n7969), .B(n12071), .Y(n8211) );
  OAI21X1 U11559 ( .A0(test_se), .A1(n12054), .B0(n7918), .Y(n8210) );
  INVX1 U11560 ( .A(n12071), .Y(n12054) );
  NOR2X1 U11561 ( .A(n11019), .B(n12072), .Y(n12071) );
  MX2X1 U11562 ( .A(n12073), .B(n12074), .S0(n7244), .Y(n12072) );
  NAND3X1 U11563 ( .A(n7575), .B(n7321), .C(n12477), .Y(n12074) );
  INVX1 U11564 ( .A(n12050), .Y(n12073) );
  NOR2X1 U11565 ( .A(n12926), .B(n12927), .Y(n12050) );
  NAND3X1 U11566 ( .A(n12932), .B(n7536), .C(n12069), .Y(n11019) );
  INVX1 U11567 ( .A(n10998), .Y(n12069) );
  NAND2X1 U11568 ( .A(n12933), .B(n12934), .Y(n10998) );
  MX2X1 U11569 ( .A(n12299), .B(g17778), .S0(n7852), .Y(n5928) );
  MX2X1 U11570 ( .A(g17722), .B(g12470), .S0(n7851), .Y(n5927) );
  MX2X1 U11571 ( .A(g12470), .B(g14828), .S0(n7851), .Y(n5926) );
  MX2X1 U11572 ( .A(g14749), .B(g17764), .S0(n7851), .Y(n5925) );
  OAI21X1 U11573 ( .A0(n12075), .A1(n12076), .B0(n12077), .Y(n5924) );
  MX2X1 U11574 ( .A(n12078), .B(n7818), .S0(n7961), .Y(n12077) );
  NAND2X1 U11575 ( .A(n12075), .B(n7424), .Y(n12078) );
  INVX1 U11576 ( .A(n12079), .Y(n12075) );
  OAI21X1 U11577 ( .A0(n7986), .A1(n7856), .B0(n12080), .Y(n5923) );
  AOI21X1 U11578 ( .A0(n12188), .A1(n7873), .B0(n12081), .Y(n12080) );
  NOR2X1 U11579 ( .A(test_se), .B(g35), .Y(n8108) );
  INVX1 U11580 ( .A(n12082), .Y(n5922) );
  AOI22X1 U11581 ( .A0(n12185), .A1(n7940), .B0(n12188), .B1(test_se), .Y(
        n12082) );
  NOR2X1 U11582 ( .A(n12083), .B(n12084), .Y(n5921) );
  MX2X1 U11583 ( .A(n12303), .B(n7424), .S0(n7961), .Y(n12084) );
  NOR2X1 U11584 ( .A(n12083), .B(n7667), .Y(n5920) );
  NOR2X1 U11585 ( .A(n12076), .B(n12079), .Y(n12083) );
  NAND4X1 U11586 ( .A(g17778), .B(g17688), .C(g14828), .D(g12470), .Y(n12079)
         );
  INVX1 U11587 ( .A(n12081), .Y(n12076) );
  NOR2X1 U11588 ( .A(n7424), .B(n7969), .Y(n12081) );
  INVX1 U11589 ( .A(n12085), .Y(n5919) );
  AOI21X1 U11590 ( .A0(n7978), .A1(n12303), .B0(n12086), .Y(n12085) );
  MX2X1 U11591 ( .A(n8249), .B(n8349), .S0(n7248), .Y(n12086) );
  INVX1 U11592 ( .A(n8252), .Y(n8349) );
  NAND2X1 U11593 ( .A(n7924), .B(n9721), .Y(n8252) );
  NOR2X1 U11594 ( .A(n9721), .B(n7963), .Y(n8249) );
  NAND2X1 U11595 ( .A(n7431), .B(n12087), .Y(n9721) );
  NAND3X1 U11596 ( .A(n12391), .B(n8615), .C(n9183), .Y(n12087) );
  INVX1 U11597 ( .A(n12088), .Y(n9183) );
  NAND4X1 U11598 ( .A(n12089), .B(n12606), .C(n12090), .D(n12608), .Y(n12088)
         );
  NOR2X1 U11599 ( .A(n12605), .B(n12610), .Y(n12090) );
  NOR2X1 U11600 ( .A(n7250), .B(n7576), .Y(n12089) );
  NOR2X1 U11601 ( .A(n7379), .B(n7247), .Y(n8615) );
  NOR2X1 U11602 ( .A(n9237), .B(test_se), .Y(n8114) );
  MX2X1 U11603 ( .A(n7248), .B(g14749), .S0(n7850), .Y(n5918) );
  INVX1 U11604 ( .A(test_se), .Y(n8104) );
  INVX1 U11605 ( .A(rst), .Y(n5917) );
  AND2X1 U11606 ( .A(n12537), .B(n12091), .Y(g34956) );
  NAND4X1 U11607 ( .A(n12539), .B(n12540), .C(n12541), .D(n7762), .Y(n12091)
         );
  AOI21X1 U11608 ( .A0(n12049), .A1(n7460), .B0(n7258), .Y(g34788) );
  INVX1 U11609 ( .A(n12092), .Y(n12049) );
  NAND3X1 U11610 ( .A(n7284), .B(n7462), .C(n12928), .Y(n12092) );
  AOI21X1 U11611 ( .A0(n12093), .A1(n12094), .B0(n12095), .Y(g34435) );
  NAND2X1 U11612 ( .A(n7384), .B(n7269), .Y(n12095) );
  NAND4X1 U11613 ( .A(n12581), .B(n9465), .C(n7236), .D(n7506), .Y(n12094) );
  NOR2X1 U11614 ( .A(n12579), .B(n12578), .Y(n9465) );
  NOR2X1 U11615 ( .A(n12576), .B(n12577), .Y(n12093) );
  INVX1 U11616 ( .A(n9987), .Y(g33959) );
  NAND2X1 U11617 ( .A(n12995), .B(n12096), .Y(n9987) );
  NAND3X1 U11618 ( .A(n13002), .B(n8632), .C(n10137), .Y(n12096) );
  INVX1 U11619 ( .A(n12097), .Y(n10137) );
  NAND4X1 U11620 ( .A(n12098), .B(n12998), .C(n12099), .D(n13000), .Y(n12097)
         );
  NOR2X1 U11621 ( .A(n12996), .B(n13001), .Y(n12099) );
  NOR2X1 U11622 ( .A(n7255), .B(n7577), .Y(n12098) );
  NOR2X1 U11623 ( .A(n7249), .B(n7380), .Y(n8632) );
  NAND2X1 U11624 ( .A(n12100), .B(n12101), .Y(g33435) );
  AOI22X1 U11625 ( .A0(n12102), .A1(n13008), .B0(n13011), .B1(n11623), .Y(
        n12101) );
  NOR2X1 U11626 ( .A(n13027), .B(n7492), .Y(n12102) );
  AOI22X1 U11627 ( .A0(n11558), .A1(n7531), .B0(n13010), .B1(n12004), .Y(
        n12100) );
  AND2X1 U11628 ( .A(n12103), .B(n12104), .Y(g33079) );
  AOI22X1 U11629 ( .A0(n12105), .A1(n13028), .B0(n11558), .B1(n7218), .Y(
        n12104) );
  NOR2X1 U11630 ( .A(n7300), .B(n7492), .Y(n11558) );
  NOR2X1 U11631 ( .A(n13018), .B(n13027), .Y(n12105) );
  AOI22X1 U11632 ( .A0(n12004), .A1(n7381), .B0(n11623), .B1(n7271), .Y(n12103) );
  NOR2X1 U11633 ( .A(n7300), .B(n13028), .Y(n11623) );
  NOR2X1 U11634 ( .A(n13028), .B(n13027), .Y(n12004) );
  NOR2X1 U11635 ( .A(n7264), .B(n10066), .Y(g32975) );
  OR2X1 U11636 ( .A(n7493), .B(n12256), .Y(n10066) );
  INVX1 U11637 ( .A(n12106), .Y(g32185) );
  NAND4X1 U11638 ( .A(n12107), .B(n12108), .C(n12109), .D(n12110), .Y(n12106)
         );
  AOI22X1 U11639 ( .A0(n12660), .A1(n12658), .B0(n12642), .B1(n12659), .Y(
        n12110) );
  AOI22X1 U11640 ( .A0(n12655), .A1(n12656), .B0(n12654), .B1(n12652), .Y(
        n12109) );
  NAND2X1 U11641 ( .A(n12643), .B(n12644), .Y(n12108) );
  AOI22X1 U11642 ( .A0(n12647), .A1(n12651), .B0(n12645), .B1(n12646), .Y(
        n12107) );
  INVX1 U11643 ( .A(n11660), .Y(g31862) );
  NAND2X1 U11644 ( .A(n12890), .B(n7421), .Y(n11660) );
  INVX1 U11645 ( .A(n12111), .Y(g31793) );
  AOI22X1 U11646 ( .A0(n8772), .A1(n12112), .B0(n12113), .B1(n8798), .Y(n12111) );
  AOI21X1 U11647 ( .A0(g35), .A1(n12670), .B0(n12114), .Y(n8798) );
  AOI22X1 U11648 ( .A0(n9975), .A1(n12115), .B0(n12116), .B1(n12117), .Y(
        n12113) );
  NAND4X1 U11649 ( .A(n12118), .B(n12119), .C(n12120), .D(n12121), .Y(n12117)
         );
  OAI21X1 U11650 ( .A0(n12679), .A1(n12678), .B0(n12677), .Y(n12120) );
  NAND2X1 U11651 ( .A(n12678), .B(n12679), .Y(n12119) );
  INVX1 U11652 ( .A(n12122), .Y(n12116) );
  INVX1 U11653 ( .A(n12118), .Y(n12115) );
  OAI21X1 U11654 ( .A0(n12670), .A1(n12123), .B0(n12114), .Y(n12112) );
  INVX1 U11655 ( .A(n8773), .Y(n12114) );
  NAND2X1 U11656 ( .A(g35), .B(n12124), .Y(n8773) );
  NAND3X1 U11657 ( .A(n7322), .B(n7620), .C(n7229), .Y(n12124) );
  AOI21X1 U11658 ( .A0(n7229), .A1(n7322), .B0(n12125), .Y(n12123) );
  AOI21X1 U11659 ( .A0(n12673), .A1(n12674), .B0(n12672), .Y(n12125) );
  INVX1 U11660 ( .A(n12126), .Y(n8772) );
  NAND3X1 U11661 ( .A(n12122), .B(n12121), .C(n12118), .Y(n12126) );
  NOR2X1 U11662 ( .A(n12675), .B(n12676), .Y(n12118) );
  INVX1 U11663 ( .A(n9975), .Y(n12121) );
  NOR2X1 U11664 ( .A(n7823), .B(n9237), .Y(n9975) );
  NAND2X1 U11665 ( .A(g35), .B(n12127), .Y(n12122) );
  NAND3X1 U11666 ( .A(n7230), .B(n7621), .C(n7331), .Y(n12127) );
  NAND3X1 U11667 ( .A(n7640), .B(n7332), .C(g35), .Y(g28042) );
  NAND3X1 U11668 ( .A(n10637), .B(n10801), .C(g35), .Y(g28041) );
  INVX1 U11669 ( .A(n8783), .Y(n10801) );
  NOR2X1 U11670 ( .A(n7689), .B(n8126), .Y(n8783) );
  NOR2X1 U11671 ( .A(n12955), .B(n12956), .Y(n8126) );
  INVX1 U11672 ( .A(n8784), .Y(n10637) );
  NOR2X1 U11673 ( .A(n7690), .B(n8132), .Y(n8784) );
  NOR2X1 U11674 ( .A(n13068), .B(n13071), .Y(n8132) );
  OAI33X1 U11675 ( .A0(n12128), .A1(n12129), .A2(n12130), .B0(n12131), .B1(
        n12132), .B2(n12133), .Y(g28030) );
  AOI21X1 U11676 ( .A0(n12134), .A1(n8800), .B0(n8801), .Y(n12132) );
  INVX1 U11677 ( .A(n12130), .Y(n8801) );
  AOI21X1 U11678 ( .A0(n12135), .A1(n12136), .B0(n12137), .Y(n12134) );
  AOI21X1 U11679 ( .A0(n7579), .A1(n7323), .B0(n12138), .Y(n12137) );
  AOI21X1 U11680 ( .A0(g35), .A1(n12136), .B0(n12135), .Y(n12138) );
  NAND2X1 U11681 ( .A(n12139), .B(n8802), .Y(n12131) );
  OAI21X1 U11682 ( .A0(n7599), .A1(n12695), .B0(n12140), .Y(n12139) );
  OR4X1 U11683 ( .A(n12136), .B(n12135), .C(n12693), .D(n12692), .Y(n12130) );
  AOI21X1 U11684 ( .A0(n7641), .A1(n12691), .B0(n9237), .Y(n12135) );
  NAND2X1 U11685 ( .A(n12690), .B(n7642), .Y(n12136) );
  AOI21X1 U11686 ( .A0(n12141), .A1(n8803), .B0(n8802), .Y(n12129) );
  NOR2X1 U11687 ( .A(n12142), .B(n12143), .Y(n8802) );
  INVX1 U11688 ( .A(n12133), .Y(n8803) );
  AOI21X1 U11689 ( .A0(n7643), .A1(n7333), .B0(n9237), .Y(n12133) );
  NAND2X1 U11690 ( .A(n12143), .B(n12142), .Y(n12141) );
  AOI21X1 U11691 ( .A0(n7644), .A1(n12689), .B0(n9237), .Y(n12142) );
  AOI21X1 U11692 ( .A0(n7645), .A1(n7334), .B0(n9237), .Y(n12143) );
  INVX1 U11693 ( .A(n8800), .Y(n12128) );
  NOR2X1 U11694 ( .A(n12140), .B(n12144), .Y(n8800) );
  AOI21X1 U11695 ( .A0(n12696), .A1(n7622), .B0(n9237), .Y(n12144) );
  AOI21X1 U11696 ( .A0(n7646), .A1(n12694), .B0(n9237), .Y(n12140) );
  INVX1 U11697 ( .A(g35), .Y(n9237) );
  AOI21X1 U11698 ( .A0(n11814), .A1(n10619), .B0(n5246), .Y(g27831) );
  INVX1 U11699 ( .A(n10587), .Y(n10619) );
  NAND2X1 U11700 ( .A(n13053), .B(n7557), .Y(n10587) );
  INVX1 U11701 ( .A(n11607), .Y(n11814) );
  NAND4X1 U11702 ( .A(n12145), .B(n13061), .C(n12146), .D(n7532), .Y(n11607)
         );
  NOR2X1 U11703 ( .A(n13016), .B(n13046), .Y(n12146) );
  NOR2X1 U11704 ( .A(n13049), .B(n7266), .Y(n12145) );
  NAND3X1 U11705 ( .A(n12147), .B(n12148), .C(g35), .Y(g26877) );
  INVX1 U11706 ( .A(n11884), .Y(n12148) );
  NOR2X1 U11707 ( .A(n12149), .B(n12150), .Y(n11884) );
  NAND4X1 U11708 ( .A(n7691), .B(n7232), .C(n7345), .D(n7208), .Y(n12150) );
  NAND4X1 U11709 ( .A(n7692), .B(n7233), .C(n7346), .D(n7209), .Y(n12149) );
  INVX1 U11710 ( .A(n11885), .Y(n12147) );
  NOR2X1 U11711 ( .A(n12151), .B(n12152), .Y(n11885) );
  NAND4X1 U11712 ( .A(n7693), .B(n7234), .C(n7347), .D(n7210), .Y(n12152) );
  NAND4X1 U11713 ( .A(n7694), .B(n7235), .C(n7348), .D(n7211), .Y(n12151) );
  NAND3X1 U11714 ( .A(n8805), .B(n8804), .C(g35), .Y(g26876) );
  OR2X1 U11715 ( .A(n12153), .B(n12154), .Y(n8804) );
  NAND4X1 U11716 ( .A(n7763), .B(n7335), .C(n7237), .D(n7212), .Y(n12154) );
  NAND4X1 U11717 ( .A(n7648), .B(n7336), .C(n7238), .D(n7213), .Y(n12153) );
  OR2X1 U11718 ( .A(n12155), .B(n12156), .Y(n8805) );
  NAND4X1 U11719 ( .A(n7337), .B(n7239), .C(n7214), .D(n7764), .Y(n12156) );
  NAND4X1 U11720 ( .A(n7649), .B(n7338), .C(n7240), .D(n7215), .Y(n12155) );
  NAND3X1 U11721 ( .A(n8807), .B(n8806), .C(g35), .Y(g26875) );
  NAND4X1 U11722 ( .A(n7765), .B(n7351), .C(n7241), .D(n7216), .Y(n8806) );
  NAND4X1 U11723 ( .A(n12797), .B(n12824), .C(n12849), .D(n12873), .Y(n8807)
         );
  NOR2X1 U11724 ( .A(n7511), .B(n12878), .Y(g25167) );
  INVX1 U11725 ( .A(n10114), .Y(g25114) );
  NAND2X1 U11726 ( .A(n12993), .B(n7366), .Y(n10114) );
  NOR2X1 U11727 ( .A(g35), .B(n7827), .Y(g21727) );
endmodule

