`timescale 1ns / 1ps

module s38584_RN320_tb;

    integer i, j, k, file;
    integer hamming_distance[11:0];
    integer hamming_weight_s38584[11:0];
    integer hamming_weight_RN320[11:0];

    reg [282:0] output_s38584[11:0];
    reg [282:0] output_RN320[11:0];

    // Inputs
    reg clk, rst, g35, g36, g6744, g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6752, g6753, test_se, test_si;

    // Outputs
    wire g7243, g7245, g7257, g7260, g7540, g7916, g7946, g8132, g8178, g8215,
        g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353, g8358, g8398,
        g8403, g8416, g8475, g8719, g8783, g8784, g8785, g8786, g8787, g8788,
        g8789, g8839, g8870, g8915, g8916, g8917, g8918, g8919, g8920, g9019,
        g9048, g9251, g9497, g9553, g9555, g9615, g9617, g9680, g9682, g9741,
        g9743, g9817, g10122, g10306, g10500, g10527, g11349, g11388, g11418,
        g11447, g11678, g11770, g12184, g12238, g12300, g12350, g12368,
        g12422, g12470, g12832, g12919, g12923, g13039, g13049, g13068,
        g13085, g13099, g13259, g13272, g13865, g13881, g13895, g13906,
        g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201,
        g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673,
        g14694, g14705, g14738, g14749, g14779, g14828, g16603, g16624,
        g16627, g16656, g16659, g16686, g16693, g16718, g16722, g16744,
        g16748, g16775, g16874, g16924, g16955, g17291, g17316, g17320,
        g17400, g17404, g17423, g17519, g17577, g17580, g17604, g17607,
        g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711,
        g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787,
        g17813, g17819, g17845, g17871, g18092, g18094, g18095, g18096,
        g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357,
        g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176,
        g21245, g21270, g21292, g21698, g21727, g23002, g23190, g23612,
        g23652, g23683, g23759, g24151, g25114, g25167, g25219, g25259,
        g25582, g25583, g25584, g25585, g25586, g25587, g25588, g25589,
        g25590, g26801, g26875, g26876, g26877, g27831, g28030, g28041,
        g28042, g28753, g29210, g29211, g29212, g29213, g29214, g29215,
        g29216, g29217, g29218, g29219, g29220, g29221, g30327, g30329,
        g30330, g30331, g30332, g31521, g31656, g31665, g31793, g31860,
        g31861, g31862, g31863, g32185, g32429, g32454, g32975, g33079,
        g33435, g33533, g33636, g33659, g33874, g33894, g33935, g33945,
        g33946, g33947, g33948, g33949, g33950, g33959, g34201, g34221,
        g34232, g34233, g34234, g34235, g34236, g34237, g34238, g34239,
        g34240, g34383, g34425, g34435, g34436, g34437, g34597, g34788,
        g34839, g34913, g34915, g34917, g34919, g34921, g34923, g34925,
        g34927, g34956, g34972;

    // Instantiate the Designs
    s38584 dut (clk, rst, g35, g36, g6744, g6745, g6746, g6747, g6748, g6749, 
        g6750, g6751, g6752, g6753, g7243, g7245, g7257, g7260, g7540, g7916, 
        g7946, g8132, g8178, g8215, g8235, g8277, g8279, g8283, g8291, g8342, 
        g8344, g8353, g8358, g8398, g8403, g8416, g8475, g8719, g8783, g8784, 
        g8785, g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916, g8917, 
        g8918, g8919, g8920, g9019, g9048, g9251, g9497, g9553, g9555, g9615, 
        g9617, g9680, g9682, g9741, g9743, g9817, g10122, g10306, g10500, 
        g10527, g11349, g11388, g11418, g11447, g11678, g11770, g12184, g12238, 
        g12300, g12350, g12368, g12422, g12470, g12832, g12919, g12923, g13039, 
        g13049, g13068, g13085, g13099, g13259, g13272, g13865, g13881, g13895, 
        g13906, g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201, 
        g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673, g14694, 
        g14705, g14738, g14749, g14779, g14828, g16603, g16624, g16627, g16656, 
        g16659, g16686, g16693, g16718, g16722, g16744, g16748, g16775, g16874, 
        g16924, g16955, g17291, g17316, g17320, g17400, g17404, g17423, g17519, 
        g17577, g17580, g17604, g17607, g17639, g17646, g17649, g17674, g17678, 
        g17685, g17688, g17711, g17715, g17722, g17739, g17743, g17760, g17764, 
        g17778, g17787, g17813, g17819, g17845, g17871, g18092, g18094, g18095, 
        g18096, g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357, 
        g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176, g21245, 
        g21270, g21292, g21698, g21727, g23002, g23190, g23612, g23652, g23683, 
        g23759, g24151, g25114, g25167, g25219, g25259, g25582, g25583, g25584, 
        g25585, g25586, g25587, g25588, g25589, g25590, g26801, g26875, g26876, 
        g26877, g27831, g28030, g28041, g28042, g28753, g29210, g29211, g29212, 
        g29213, g29214, g29215, g29216, g29217, g29218, g29219, g29220, g29221, 
        g30327, g30329, g30330, g30331, g30332, g31521, g31656, g31665, g31793, 
        g31860, g31861, g31862, g31863, g32185, g32429, g32454, g32975, g33079, 
        g33435, g33533, g33636, g33659, g33874, g33894, g33935, g33945, g33946, 
        g33947, g33948, g33949, g33950, g33959, g34201, g34221, g34232, g34233, 
        g34234, g34235, g34236, g34237, g34238, g34239, g34240, g34383, g34425, 
        g34435, g34436, g34437, g34597, g34788, g34839, g34913, g34915, g34917, 
        g34919, g34921, g34923, g34925, g34927, g34956, g34972, test_se, 
        test_si );


    // Inputs
    reg g35_RN, g36_RN, g6744_RN, g6745_RN, g6746_RN, g6747_RN, g6748_RN, g6749_RN, g6750_RN, g6751_RN, g6752_RN, g6753_RN, test_se_RN, test_si_RN;
    reg [0:31] keyinput;
    // Outputs
    wire g7243_RN, g7245_RN, g7257_RN, g7260_RN, g7540_RN, g7916_RN, g7946_RN, g8132_RN, g8178_RN, g8215_RN,
        g8235_RN, g8277_RN, g8279_RN, g8283_RN, g8291_RN, g8342_RN, g8344_RN, g8353_RN, g8358_RN, g8398_RN,
        g8403_RN, g8416_RN, g8475_RN, g8719_RN, g8783_RN, g8784_RN, g8785_RN, g8786_RN, g8787_RN, g8788_RN,
        g8789_RN, g8839_RN, g8870_RN, g8915_RN, g8916_RN, g8917_RN, g8918_RN, g8919_RN, g8920_RN, g9019_RN,
        g9048_RN, g9251_RN, g9497_RN, g9553_RN, g9555_RN, g9615_RN, g9617_RN, g9680_RN, g9682_RN, g9741_RN,
        g9743_RN, g9817_RN, g10122_RN, g10306_RN, g10500_RN, g10527_RN, g11349_RN, g11388_RN, g11418_RN,
        g11447_RN, g11678_RN, g11770_RN, g12184_RN, g12238_RN, g12300_RN, g12350_RN, g12368_RN,
        g12422_RN, g12470_RN, g12832_RN, g12919_RN, g12923_RN, g13039_RN, g13049_RN, g13068_RN,
        g13085_RN, g13099_RN, g13259_RN, g13272_RN, g13865_RN, g13881_RN, g13895_RN, g13906_RN,
        g13926_RN, g13966_RN, g14096_RN, g14125_RN, g14147_RN, g14167_RN, g14189_RN, g14201_RN,
        g14217_RN, g14421_RN, g14451_RN, g14518_RN, g14597_RN, g14635_RN, g14662_RN, g14673_RN,
        g14694_RN, g14705_RN, g14738_RN, g14749_RN, g14779_RN, g14828_RN, g16603_RN, g16624_RN,
        g16627_RN, g16656_RN, g16659_RN, g16686_RN, g16693_RN, g16718_RN, g16722_RN, g16744_RN,
        g16748_RN, g16775_RN, g16874_RN, g16924_RN, g16955_RN, g17291_RN, g17316_RN, g17320_RN,
        g17400_RN, g17404_RN, g17423_RN, g17519_RN, g17577_RN, g17580_RN, g17604_RN, g17607_RN,
        g17639_RN, g17646_RN, g17649_RN, g17674_RN, g17678_RN, g17685_RN, g17688_RN, g17711_RN,
        g17715_RN, g17722_RN, g17739_RN, g17743_RN, g17760_RN, g17764_RN, g17778_RN, g17787_RN,
        g17813_RN, g17819_RN, g17845_RN, g17871_RN, g18092_RN, g18094_RN, g18095_RN, g18096_RN,
        g18097_RN, g18098_RN, g18099_RN, g18100_RN, g18101_RN, g18881_RN, g19334_RN, g19357_RN,
        g20049_RN, g20557_RN, g20652_RN, g20654_RN, g20763_RN, g20899_RN, g20901_RN, g21176_RN,
        g21245_RN, g21270_RN, g21292_RN, g21698_RN, g21727_RN, g23002_RN, g23190_RN, g23612_RN,
        g23652_RN, g23683_RN, g23759_RN, g24151_RN, g25114_RN, g25167_RN, g25219_RN, g25259_RN,
        g25582_RN, g25583_RN, g25584_RN, g25585_RN, g25586_RN, g25587_RN, g25588_RN, g25589_RN,
        g25590_RN, g26801_RN, g26875_RN, g26876_RN, g26877_RN, g27831_RN, g28030_RN, g28041_RN,
        g28042_RN, g28753_RN, g29210_RN, g29211_RN, g29212_RN, g29213_RN, g29214_RN, g29215_RN,
        g29216_RN, g29217_RN, g29218_RN, g29219_RN, g29220_RN, g29221_RN, g30327_RN, g30329_RN,
        g30330_RN, g30331_RN, g30332_RN, g31521_RN, g31656_RN, g31665_RN, g31793_RN, g31860_RN,
        g31861_RN, g31862_RN, g31863_RN, g32185_RN, g32429_RN, g32454_RN, g32975_RN, g33079_RN,
        g33435_RN, g33533_RN, g33636_RN, g33659_RN, g33874_RN, g33894_RN, g33935_RN, g33945_RN,
        g33946_RN, g33947_RN, g33948_RN, g33949_RN, g33950_RN, g33959_RN, g34201_RN, g34221_RN,
        g34232_RN, g34233_RN, g34234_RN, g34235_RN, g34236_RN, g34237_RN, g34238_RN, g34239_RN,
        g34240_RN, g34383_RN, g34425_RN, g34435_RN, g34436_RN, g34437_RN, g34597_RN, g34788_RN,
        g34839_RN, g34913_RN, g34915_RN, g34917_RN, g34919_RN, g34921_RN, g34923_RN, g34925_RN,
        g34927_RN, g34956_RN, g34972_RN;


    s38584_RN320 dut_RN (clk, rst, g35_RN, g36_RN, g6744_RN, g6745_RN, g6746_RN, g6747_RN, g6748_RN, g6749_RN,
        g6750_RN, g6751_RN, g6752_RN, g6753_RN, g7243_RN, g7245_RN, g7257_RN, g7260_RN, g7540_RN, g7916_RN, 
        g7946_RN, g8132_RN, g8178_RN, g8215_RN, g8235_RN, g8277_RN, g8279_RN, g8283_RN, g8291_RN, g8342_RN, 
        g8344_RN, g8353_RN, g8358_RN, g8398_RN, g8403_RN, g8416_RN, g8475_RN, g8719_RN, g8783_RN, g8784_RN, 
        g8785_RN, g8786_RN, g8787_RN, g8788_RN, g8789_RN, g8839_RN, g8870_RN, g8915_RN, g8916_RN, g8917_RN, 
        g8918_RN, g8919_RN, g8920_RN, g9019_RN, g9048_RN, g9251_RN, g9497_RN, g9553_RN, g9555_RN, g9615_RN, 
        g9617_RN, g9680_RN, g9682_RN, g9741_RN, g9743_RN, g9817_RN, g10122_RN, g10306_RN, g10500_RN, 
        g10527_RN, g11349_RN, g11388_RN, g11418_RN, g11447_RN, g11678_RN, g11770_RN, g12184_RN, g12238_RN, 
        g12300_RN, g12350_RN, g12368_RN, g12422_RN, g12470_RN, g12832_RN, g12919_RN, g12923_RN, g13039_RN, 
        g13049_RN, g13068_RN, g13085_RN, g13099_RN, g13259_RN, g13272_RN, g13865_RN, g13881_RN, g13895_RN, 
        g13906_RN, g13926_RN, g13966_RN, g14096_RN, g14125_RN, g14147_RN, g14167_RN, g14189_RN, g14201_RN, 
        g14217_RN, g14421_RN, g14451_RN, g14518_RN, g14597_RN, g14635_RN, g14662_RN, g14673_RN, g14694_RN, 
        g14705_RN, g14738_RN, g14749_RN, g14779_RN, g14828_RN, g16603_RN, g16624_RN, g16627_RN, g16656_RN, 
        g16659_RN, g16686_RN, g16693_RN, g16718_RN, g16722_RN, g16744_RN, g16748_RN, g16775_RN, g16874_RN, 
        g16924_RN, g16955_RN, g17291_RN, g17316_RN, g17320_RN, g17400_RN, g17404_RN, g17423_RN, g17519_RN, 
        g17577_RN, g17580_RN, g17604_RN, g17607_RN, g17639_RN, g17646_RN, g17649_RN, g17674_RN, g17678_RN, 
        g17685_RN, g17688_RN, g17711_RN, g17715_RN, g17722_RN, g17739_RN, g17743_RN, g17760_RN, g17764_RN, 
        g17778_RN, g17787_RN, g17813_RN, g17819_RN, g17845_RN, g17871_RN, g18092_RN, g18094_RN, g18095_RN, 
        g18096_RN, g18097_RN, g18098_RN, g18099_RN, g18100_RN, g18101_RN, g18881_RN, g19334_RN, g19357_RN, 
        g20049_RN, g20557_RN, g20652_RN, g20654_RN, g20763_RN, g20899_RN, g20901_RN, g21176_RN, g21245_RN, 
        g21270_RN, g21292_RN, g21698_RN, g21727_RN, g23002_RN, g23190_RN, g23612_RN, g23652_RN, g23683_RN, 
        g23759_RN, g24151_RN, g25114_RN, g25167_RN, g25219_RN, g25259_RN, g25582_RN, g25583_RN, g25584_RN, 
        g25585_RN, g25586_RN, g25587_RN, g25588_RN, g25589_RN, g25590_RN, g26801_RN, g26875_RN, g26876_RN, 
        g26877_RN, g27831_RN, g28030_RN, g28041_RN, g28042_RN, g28753_RN, g29210_RN, g29211_RN, g29212_RN, 
        g29213_RN, g29214_RN, g29215_RN, g29216_RN, g29217_RN, g29218_RN, g29219_RN, g29220_RN, g29221_RN, 
        g30327_RN, g30329_RN, g30330_RN, g30331_RN, g30332_RN, g31521_RN, g31656_RN, g31665_RN, g31793_RN, 
        g31860_RN, g31861_RN, g31862_RN, g31863_RN, g32185_RN, g32429_RN, g32454_RN, g32975_RN, g33079_RN, 
        g33435_RN, g33533_RN, g33636_RN, g33659_RN, g33874_RN, g33894_RN, g33935_RN, g33945_RN, g33946_RN, 
        g33947_RN, g33948_RN, g33949_RN, g33950_RN, g33959_RN, g34201_RN, g34221_RN, g34232_RN, g34233_RN, 
        g34234_RN, g34235_RN, g34236_RN, g34237_RN, g34238_RN, g34239_RN, g34240_RN, g34383_RN, g34425_RN, 
        g34435_RN, g34436_RN, g34437_RN, g34597_RN, g34788_RN, g34839_RN, g34913_RN, g34915_RN, g34917_RN, 
        g34919_RN, g34921_RN, g34923_RN, g34925_RN, g34927_RN, g34956_RN, g34972_RN, test_se_RN, 
        test_si_RN , keyinput);

    always // clock with period 1000ns
    begin
        clk = 1;
        #500;
        clk = !clk;
        #500;
    end
    
    // Test Patterns
    initial 
    begin

        // Create a file for writing the outputs of the testbench
        file = $fopen("tb_s38584-RN320.txt", "w");

        // Flash the reset on the DUT
        rst = 1;
        #1000;
        rst = 0;
        
        for (j=0; j < 12; j = j+1)
        begin

            // initialize all the distance and weights to zero
            hamming_distance[j] = 0;
            hamming_weight_s38584[j] = 0;
            hamming_weight_RN320[j] = 0;

        end

        for (i=0; i < 12; i = i+1)
        begin

            // Have the first test be non random.
            if (i < 2)

                // First index, test all ones
                if (i==0)
                begin

                    // assign all 1's to the inputs
                    g35 = 1;
                    g36 = 1;
                    g6744 = 1;
                    g6745 = 1;
                    g6746 = 1;
                    g6747 = 1;
                    g6748 = 1;
                    g6749 = 1;
                    g6750 = 1;
                    g6751 = 1;
                    g6752 = 1;
                    g6753 = 1;
                    test_se = 1;
                    test_si = 1;

                    g35_RN = 1;
                    g36_RN = 1;
                    g6744_RN = 1;
                    g6745_RN = 1;
                    g6746_RN = 1;
                    g6747_RN = 1;
                    g6748_RN = 1;
                    g6749_RN = 1;
                    g6750_RN = 1;
                    g6751_RN = 1;
                    g6752_RN = 1;
                    g6753_RN = 1;
                    test_se_RN = 1;
                    test_si_RN = 1;
                    keyinput = 32'hffffffff';
                end

                // Second index, test all zeros
                else
                begin

                    // assign all 0's to the inputs
                    g35 = 0;
                    g36 = 0;
                    g6744 = 0;
                    g6745 = 0;
                    g6746 = 0;
                    g6747 = 0;
                    g6748 = 0;
                    g6749 = 0;
                    g6750 = 0;
                    g6751 = 0;
                    g6752 = 0;
                    g6753 = 0;
                    test_se = 0; 
                    test_si = 0;

                    g35_RN = 0;
                    g36_RN = 0;
                    g6744_RN = 0;
                    g6745_RN = 0;
                    g6746_RN = 0;
                    g6747_RN = 0;
                    g6748_RN = 0;
                    g6749_RN = 0;
                    g6750_RN = 0;
                    g6751_RN = 0;
                    g6752_RN = 0;
                    g6753_RN = 0;
                    test_se_RN = 0;
                    test_si_RN = 0;
                    keyinput = 32'h00000000';

                end

            else
            begin
                // assign random data
                {g35, g36, g6744, g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6752, g6753, test_se, test_si} = $random;
                                    
                    // assign the same data to the RN inputs
                    g35_RN = g35;
                    g36_RN = g36;
                    g6744_RN = g6744;
                    g6745_RN = g6745;
                    g6746_RN = g6746;
                    g6747_RN = g6747;
                    g6748_RN = g6748;
                    g6749_RN = g6749;
                    g6750_RN = g6750;
                    g6751_RN = g6751;
                    g6752_RN = g6752;
                    g6753_RN = g6753;
                    test_se_RN = test_se;
                    test_si_RN = test_si;
                    keyinput = $random;

            end
            
            // write to the file 
            $fwrite(file,"Input Pattern s38584: %b\n", {g35, g36, g6744, g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6752, g6753, test_se, test_si});
            $fwrite(file,"Output Pattern s38584: %b\n", {g7243, g7245, g7257, g7260, g7540, g7916, g7946, g8132, g8178, g8215,
                                                    g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353, g8358, g8398,
                                                    g8403, g8416, g8475, g8719, g8783, g8784, g8785, g8786, g8787, g8788,
                                                    g8789, g8839, g8870, g8915, g8916, g8917, g8918, g8919, g8920, g9019,
                                                    g9048, g9251, g9497, g9553, g9555, g9615, g9617, g9680, g9682, g9741,
                                                    g9743, g9817, g10122, g10306, g10500, g10527, g11349, g11388, g11418,
                                                    g11447, g11678, g11770, g12184, g12238, g12300, g12350, g12368,
                                                    g12422, g12470, g12832, g12919, g12923, g13039, g13049, g13068,
                                                    g13085, g13099, g13259, g13272, g13865, g13881, g13895, g13906,
                                                    g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201,
                                                    g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673,
                                                    g14694, g14705, g14738, g14749, g14779, g14828, g16603, g16624,
                                                    g16627, g16656, g16659, g16686, g16693, g16718, g16722, g16744,
                                                    g16748, g16775, g16874, g16924, g16955, g17291, g17316, g17320,
                                                    g17400, g17404, g17423, g17519, g17577, g17580, g17604, g17607,
                                                    g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711,
                                                    g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787,
                                                    g17813, g17819, g17845, g17871, g18092, g18094, g18095, g18096,
                                                    g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357,
                                                    g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176,
                                                    g21245, g21270, g21292, g21698, g21727, g23002, g23190, g23612,
                                                    g23652, g23683, g23759, g24151, g25114, g25167, g25219, g25259,
                                                    g25582, g25583, g25584, g25585, g25586, g25587, g25588, g25589,
                                                    g25590, g26801, g26875, g26876, g26877, g27831, g28030, g28041,
                                                    g28042, g28753, g29210, g29211, g29212, g29213, g29214, g29215,
                                                    g29216, g29217, g29218, g29219, g29220, g29221, g30327, g30329,
                                                    g30330, g30331, g30332, g31521, g31656, g31665, g31793, g31860,
                                                    g31861, g31862, g31863, g32185, g32429, g32454, g32975, g33079,
                                                    g33435, g33533, g33636, g33659, g33874, g33894, g33935, g33945,
                                                    g33946, g33947, g33948, g33949, g33950, g33959, g34201, g34221,
                                                    g34232, g34233, g34234, g34235, g34236, g34237, g34238, g34239,
                                                    g34240, g34383, g34425, g34435, g34436, g34437, g34597, g34788,
                                                    g34839, g34913, g34915, g34917, g34919, g34921, g34923, g34925,
                                                    g34927, g34956, g34972});

            $fwrite(file,"Input Pattern RN320: %b\n", {g35_RN, g36_RN, g6744_RN, g6745_RN, g6746_RN, g6747_RN, g6748_RN, g6749_RN, g6750_RN, g6751_RN, g6752_RN, g6753_RN, test_se_RN, test_si_RN, keyinput});
            $fwrite(file,"Output Pattern RN320: %b\n", {g7243_RN, g7245_RN, g7257_RN, g7260_RN, g7540_RN, g7916_RN, g7946_RN, g8132_RN, g8178_RN, g8215_RN,
                                                        g8235_RN, g8277_RN, g8279_RN, g8283_RN, g8291_RN, g8342_RN, g8344_RN, g8353_RN, g8358_RN, g8398_RN,
                                                        g8403_RN, g8416_RN, g8475_RN, g8719_RN, g8783_RN, g8784_RN, g8785_RN, g8786_RN, g8787_RN, g8788_RN,
                                                        g8789_RN, g8839_RN, g8870_RN, g8915_RN, g8916_RN, g8917_RN, g8918_RN, g8919_RN, g8920_RN, g9019_RN,
                                                        g9048_RN, g9251_RN, g9497_RN, g9553_RN, g9555_RN, g9615_RN, g9617_RN, g9680_RN, g9682_RN, g9741_RN,
                                                        g9743_RN, g9817_RN, g10122_RN, g10306_RN, g10500_RN, g10527_RN, g11349_RN, g11388_RN, g11418_RN,
                                                        g11447_RN, g11678_RN, g11770_RN, g12184_RN, g12238_RN, g12300_RN, g12350_RN, g12368_RN,
                                                        g12422_RN, g12470_RN, g12832_RN, g12919_RN, g12923_RN, g13039_RN, g13049_RN, g13068_RN,
                                                        g13085_RN, g13099_RN, g13259_RN, g13272_RN, g13865_RN, g13881_RN, g13895_RN, g13906_RN,
                                                        g13926_RN, g13966_RN, g14096_RN, g14125_RN, g14147_RN, g14167_RN, g14189_RN, g14201_RN,
                                                        g14217_RN, g14421_RN, g14451_RN, g14518_RN, g14597_RN, g14635_RN, g14662_RN, g14673_RN,
                                                        g14694_RN, g14705_RN, g14738_RN, g14749_RN, g14779_RN, g14828_RN, g16603_RN, g16624_RN,
                                                        g16627_RN, g16656_RN, g16659_RN, g16686_RN, g16693_RN, g16718_RN, g16722_RN, g16744_RN,
                                                        g16748_RN, g16775_RN, g16874_RN, g16924_RN, g16955_RN, g17291_RN, g17316_RN, g17320_RN,
                                                        g17400_RN, g17404_RN, g17423_RN, g17519_RN, g17577_RN, g17580_RN, g17604_RN, g17607_RN,
                                                        g17639_RN, g17646_RN, g17649_RN, g17674_RN, g17678_RN, g17685_RN, g17688_RN, g17711_RN,
                                                        g17715_RN, g17722_RN, g17739_RN, g17743_RN, g17760_RN, g17764_RN, g17778_RN, g17787_RN,
                                                        g17813_RN, g17819_RN, g17845_RN, g17871_RN, g18092_RN, g18094_RN, g18095_RN, g18096_RN,
                                                        g18097_RN, g18098_RN, g18099_RN, g18100_RN, g18101_RN, g18881_RN, g19334_RN, g19357_RN,
                                                        g20049_RN, g20557_RN, g20652_RN, g20654_RN, g20763_RN, g20899_RN, g20901_RN, g21176_RN,
                                                        g21245_RN, g21270_RN, g21292_RN, g21698_RN, g21727_RN, g23002_RN, g23190_RN, g23612_RN,
                                                        g23652_RN, g23683_RN, g23759_RN, g24151_RN, g25114_RN, g25167_RN, g25219_RN, g25259_RN,
                                                        g25582_RN, g25583_RN, g25584_RN, g25585_RN, g25586_RN, g25587_RN, g25588_RN, g25589_RN,
                                                        g25590_RN, g26801_RN, g26875_RN, g26876_RN, g26877_RN, g27831_RN, g28030_RN, g28041_RN,
                                                        g28042_RN, g28753_RN, g29210_RN, g29211_RN, g29212_RN, g29213_RN, g29214_RN, g29215_RN,
                                                        g29216_RN, g29217_RN, g29218_RN, g29219_RN, g29220_RN, g29221_RN, g30327_RN, g30329_RN,
                                                        g30330_RN, g30331_RN, g30332_RN, g31521_RN, g31656_RN, g31665_RN, g31793_RN, g31860_RN,
                                                        g31861_RN, g31862_RN, g31863_RN, g32185_RN, g32429_RN, g32454_RN, g32975_RN, g33079_RN,
                                                        g33435_RN, g33533_RN, g33636_RN, g33659_RN, g33874_RN, g33894_RN, g33935_RN, g33945_RN,
                                                        g33946_RN, g33947_RN, g33948_RN, g33949_RN, g33950_RN, g33959_RN, g34201_RN, g34221_RN,
                                                        g34232_RN, g34233_RN, g34234_RN, g34235_RN, g34236_RN, g34237_RN, g34238_RN, g34239_RN,
                                                        g34240_RN, g34383_RN, g34425_RN, g34435_RN, g34436_RN, g34437_RN, g34597_RN, g34788_RN,
                                                        g34839_RN, g34913_RN, g34915_RN, g34917_RN, g34919_RN, g34921_RN, g34923_RN, g34925_RN,
                                                        g34927_RN, g34956_RN, g34972_RN});




            output_s38584[i] = {g7243, g7245, g7257, g7260, g7540, g7916, g7946, g8132, g8178, g8215,
                                g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353, g8358, g8398,
                                g8403, g8416, g8475, g8719, g8783, g8784, g8785, g8786, g8787, g8788,
                                g8789, g8839, g8870, g8915, g8916, g8917, g8918, g8919, g8920, g9019,
                                g9048, g9251, g9497, g9553, g9555, g9615, g9617, g9680, g9682, g9741,
                                g9743, g9817, g10122, g10306, g10500, g10527, g11349, g11388, g11418,
                                g11447, g11678, g11770, g12184, g12238, g12300, g12350, g12368,
                                g12422, g12470, g12832, g12919, g12923, g13039, g13049, g13068,
                                g13085, g13099, g13259, g13272, g13865, g13881, g13895, g13906,
                                g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201,
                                g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673,
                                g14694, g14705, g14738, g14749, g14779, g14828, g16603, g16624,
                                g16627, g16656, g16659, g16686, g16693, g16718, g16722, g16744,
                                g16748, g16775, g16874, g16924, g16955, g17291, g17316, g17320,
                                g17400, g17404, g17423, g17519, g17577, g17580, g17604, g17607,
                                g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711,
                                g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787,
                                g17813, g17819, g17845, g17871, g18092, g18094, g18095, g18096,
                                g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357,
                                g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176,
                                g21245, g21270, g21292, g21698, g21727, g23002, g23190, g23612,
                                g23652, g23683, g23759, g24151, g25114, g25167, g25219, g25259,
                                g25582, g25583, g25584, g25585, g25586, g25587, g25588, g25589,
                                g25590, g26801, g26875, g26876, g26877, g27831, g28030, g28041,
                                g28042, g28753, g29210, g29211, g29212, g29213, g29214, g29215,
                                g29216, g29217, g29218, g29219, g29220, g29221, g30327, g30329,
                                g30330, g30331, g30332, g31521, g31656, g31665, g31793, g31860,
                                g31861, g31862, g31863, g32185, g32429, g32454, g32975, g33079,
                                g33435, g33533, g33636, g33659, g33874, g33894, g33935, g33945,
                                g33946, g33947, g33948, g33949, g33950, g33959, g34201, g34221,
                                g34232, g34233, g34234, g34235, g34236, g34237, g34238, g34239,
                                g34240, g34383, g34425, g34435, g34436, g34437, g34597, g34788,
                                g34839, g34913, g34915, g34917, g34919, g34921, g34923, g34925,
                                g34927, g34956, g34972};

            output_RN320[i] = g7243_RN, g7245_RN, g7257_RN, g7260_RN, g7540_RN, g7916_RN, g7946_RN, g8132_RN, g8178_RN, g8215_RN,
                                g8235_RN, g8277_RN, g8279_RN, g8283_RN, g8291_RN, g8342_RN, g8344_RN, g8353_RN, g8358_RN, g8398_RN,
                                g8403_RN, g8416_RN, g8475_RN, g8719_RN, g8783_RN, g8784_RN, g8785_RN, g8786_RN, g8787_RN, g8788_RN,
                                g8789_RN, g8839_RN, g8870_RN, g8915_RN, g8916_RN, g8917_RN, g8918_RN, g8919_RN, g8920_RN, g9019_RN,
                                g9048_RN, g9251_RN, g9497_RN, g9553_RN, g9555_RN, g9615_RN, g9617_RN, g9680_RN, g9682_RN, g9741_RN,
                                g9743_RN, g9817_RN, g10122_RN, g10306_RN, g10500_RN, g10527_RN, g11349_RN, g11388_RN, g11418_RN,
                                g11447_RN, g11678_RN, g11770_RN, g12184_RN, g12238_RN, g12300_RN, g12350_RN, g12368_RN,
                                g12422_RN, g12470_RN, g12832_RN, g12919_RN, g12923_RN, g13039_RN, g13049_RN, g13068_RN,
                                g13085_RN, g13099_RN, g13259_RN, g13272_RN, g13865_RN, g13881_RN, g13895_RN, g13906_RN,
                                g13926_RN, g13966_RN, g14096_RN, g14125_RN, g14147_RN, g14167_RN, g14189_RN, g14201_RN,
                                g14217_RN, g14421_RN, g14451_RN, g14518_RN, g14597_RN, g14635_RN, g14662_RN, g14673_RN,
                                g14694_RN, g14705_RN, g14738_RN, g14749_RN, g14779_RN, g14828_RN, g16603_RN, g16624_RN,
                                g16627_RN, g16656_RN, g16659_RN, g16686_RN, g16693_RN, g16718_RN, g16722_RN, g16744_RN,
                                g16748_RN, g16775_RN, g16874_RN, g16924_RN, g16955_RN, g17291_RN, g17316_RN, g17320_RN,
                                g17400_RN, g17404_RN, g17423_RN, g17519_RN, g17577_RN, g17580_RN, g17604_RN, g17607_RN,
                                g17639_RN, g17646_RN, g17649_RN, g17674_RN, g17678_RN, g17685_RN, g17688_RN, g17711_RN,
                                g17715_RN, g17722_RN, g17739_RN, g17743_RN, g17760_RN, g17764_RN, g17778_RN, g17787_RN,
                                g17813_RN, g17819_RN, g17845_RN, g17871_RN, g18092_RN, g18094_RN, g18095_RN, g18096_RN,
                                g18097_RN, g18098_RN, g18099_RN, g18100_RN, g18101_RN, g18881_RN, g19334_RN, g19357_RN,
                                g20049_RN, g20557_RN, g20652_RN, g20654_RN, g20763_RN, g20899_RN, g20901_RN, g21176_RN,
                                g21245_RN, g21270_RN, g21292_RN, g21698_RN, g21727_RN, g23002_RN, g23190_RN, g23612_RN,
                                g23652_RN, g23683_RN, g23759_RN, g24151_RN, g25114_RN, g25167_RN, g25219_RN, g25259_RN,
                                g25582_RN, g25583_RN, g25584_RN, g25585_RN, g25586_RN, g25587_RN, g25588_RN, g25589_RN,
                                g25590_RN, g26801_RN, g26875_RN, g26876_RN, g26877_RN, g27831_RN, g28030_RN, g28041_RN,
                                g28042_RN, g28753_RN, g29210_RN, g29211_RN, g29212_RN, g29213_RN, g29214_RN, g29215_RN,
                                g29216_RN, g29217_RN, g29218_RN, g29219_RN, g29220_RN, g29221_RN, g30327_RN, g30329_RN,
                                g30330_RN, g30331_RN, g30332_RN, g31521_RN, g31656_RN, g31665_RN, g31793_RN, g31860_RN,
                                g31861_RN, g31862_RN, g31863_RN, g32185_RN, g32429_RN, g32454_RN, g32975_RN, g33079_RN,
                                g33435_RN, g33533_RN, g33636_RN, g33659_RN, g33874_RN, g33894_RN, g33935_RN, g33945_RN,
                                g33946_RN, g33947_RN, g33948_RN, g33949_RN, g33950_RN, g33959_RN, g34201_RN, g34221_RN,
                                g34232_RN, g34233_RN, g34234_RN, g34235_RN, g34236_RN, g34237_RN, g34238_RN, g34239_RN,
                                g34240_RN, g34383_RN, g34425_RN, g34435_RN, g34436_RN, g34437_RN, g34597_RN, g34788_RN,
                                g34839_RN, g34913_RN, g34915_RN, g34917_RN, g34919_RN, g34921_RN, g34923_RN, g34925_RN,
                                g34927_RN, g34956_RN, g34972_RN};

            // calculate the hamming weight of output of s38584
            for (k=0; K < 283; k = k+1)
            begin
                
                // if the output is equal to one, increase the weight
                if (output_s38584[i][k] == 1'b1)
                begin
                    hamming_weight_s38584[i] = hamming_weight_s38584[i] + 1;
                end

            end
            
            // calculate the hamming weight of output of RN320
            for (k=0; K < 283; k = k+1)
            begin
                
                // if the output is equal to one, increase the weight
                if (output_RN320[i][k] == 1'b1)
                begin
                    hamming_weight_RN320[i] = hamming_weight_RN320[i] + 1;
                end
                
            end

            // calculate the hamming distance between s38584 and RN320
            for (k=0; K < 283; k = k+1)
            begin
                
                // if the exclusive OR of the two outputs is equal to one, increase the distance
                if ( (output_RN320[i][k] ^ output_s38584[i][k])  == 1'b1)
                begin
                    hamming_distance[i] = hamming_distance[i] + 1;
                end
        
            end

            $display("Hamming Weight S38584[%d]: %d\n", i, hamming_weight_s38584[i]);
            $display("Hamming Weight RN320[%d]: %d\n", i, hamming_weight_RN320[i]);
            $display("Hamming Dsitance[%d]: %d\n", i, hamming_distance[i]);

            $fwrite(file, "Hamming Weight S38584[%d]: %d\n", i, hamming_weight_s38584[i]);
            $fwrite(file, "Hamming Weight RN320[%d]: %d\n", i, hamming_weight_RN320[i]);
            $fwrite(file, "Hamming Dsitance[%d]: %d\n", i, hamming_distance[i]);
        
            // wait 5000 ns before the next iteration
            #5000;

        end    

    // Close the file
    $fclose(file);
    $finish;
    end

endmodule