`timescale 1ns / 1ps

module s38584_tb;

    integer i, file;

    // Inputs
    reg clk, rst, g35, g36, g6744, g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6752, g6753, test_se, test_si;

    // Outputs
    wire g7243, g7245, g7257, g7260, g7540, g7916, g7946, g8132, g8178, g8215,
        g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353, g8358, g8398,
        g8403, g8416, g8475, g8719, g8783, g8784, g8785, g8786, g8787, g8788,
        g8789, g8839, g8870, g8915, g8916, g8917, g8918, g8919, g8920, g9019,
        g9048, g9251, g9497, g9553, g9555, g9615, g9617, g9680, g9682, g9741,
        g9743, g9817, g10122, g10306, g10500, g10527, g11349, g11388, g11418,
        g11447, g11678, g11770, g12184, g12238, g12300, g12350, g12368,
        g12422, g12470, g12832, g12919, g12923, g13039, g13049, g13068,
        g13085, g13099, g13259, g13272, g13865, g13881, g13895, g13906,
        g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201,
        g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673,
        g14694, g14705, g14738, g14749, g14779, g14828, g16603, g16624,
        g16627, g16656, g16659, g16686, g16693, g16718, g16722, g16744,
        g16748, g16775, g16874, g16924, g16955, g17291, g17316, g17320,
        g17400, g17404, g17423, g17519, g17577, g17580, g17604, g17607,
        g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711,
        g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787,
        g17813, g17819, g17845, g17871, g18092, g18094, g18095, g18096,
        g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357,
        g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176,
        g21245, g21270, g21292, g21698, g21727, g23002, g23190, g23612,
        g23652, g23683, g23759, g24151, g25114, g25167, g25219, g25259,
        g25582, g25583, g25584, g25585, g25586, g25587, g25588, g25589,
        g25590, g26801, g26875, g26876, g26877, g27831, g28030, g28041,
        g28042, g28753, g29210, g29211, g29212, g29213, g29214, g29215,
        g29216, g29217, g29218, g29219, g29220, g29221, g30327, g30329,
        g30330, g30331, g30332, g31521, g31656, g31665, g31793, g31860,
        g31861, g31862, g31863, g32185, g32429, g32454, g32975, g33079,
        g33435, g33533, g33636, g33659, g33874, g33894, g33935, g33945,
        g33946, g33947, g33948, g33949, g33950, g33959, g34201, g34221,
        g34232, g34233, g34234, g34235, g34236, g34237, g34238, g34239,
        g34240, g34383, g34425, g34435, g34436, g34437, g34597, g34788,
        g34839, g34913, g34915, g34917, g34919, g34921, g34923, g34925,
        g34927, g34956, g34972;

    // Instantiate the Design
    s38584 dut (clk, rst, g35, g36, g6744, g6745, g6746, g6747, g6748, g6749, 
        g6750, g6751, g6752, g6753, g7243, g7245, g7257, g7260, g7540, g7916, 
        g7946, g8132, g8178, g8215, g8235, g8277, g8279, g8283, g8291, g8342, 
        g8344, g8353, g8358, g8398, g8403, g8416, g8475, g8719, g8783, g8784, 
        g8785, g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916, g8917, 
        g8918, g8919, g8920, g9019, g9048, g9251, g9497, g9553, g9555, g9615, 
        g9617, g9680, g9682, g9741, g9743, g9817, g10122, g10306, g10500, 
        g10527, g11349, g11388, g11418, g11447, g11678, g11770, g12184, g12238, 
        g12300, g12350, g12368, g12422, g12470, g12832, g12919, g12923, g13039, 
        g13049, g13068, g13085, g13099, g13259, g13272, g13865, g13881, g13895, 
        g13906, g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201, 
        g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673, g14694, 
        g14705, g14738, g14749, g14779, g14828, g16603, g16624, g16627, g16656, 
        g16659, g16686, g16693, g16718, g16722, g16744, g16748, g16775, g16874, 
        g16924, g16955, g17291, g17316, g17320, g17400, g17404, g17423, g17519, 
        g17577, g17580, g17604, g17607, g17639, g17646, g17649, g17674, g17678, 
        g17685, g17688, g17711, g17715, g17722, g17739, g17743, g17760, g17764, 
        g17778, g17787, g17813, g17819, g17845, g17871, g18092, g18094, g18095, 
        g18096, g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357, 
        g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176, g21245, 
        g21270, g21292, g21698, g21727, g23002, g23190, g23612, g23652, g23683, 
        g23759, g24151, g25114, g25167, g25219, g25259, g25582, g25583, g25584, 
        g25585, g25586, g25587, g25588, g25589, g25590, g26801, g26875, g26876, 
        g26877, g27831, g28030, g28041, g28042, g28753, g29210, g29211, g29212, 
        g29213, g29214, g29215, g29216, g29217, g29218, g29219, g29220, g29221, 
        g30327, g30329, g30330, g30331, g30332, g31521, g31656, g31665, g31793, 
        g31860, g31861, g31862, g31863, g32185, g32429, g32454, g32975, g33079, 
        g33435, g33533, g33636, g33659, g33874, g33894, g33935, g33945, g33946, 
        g33947, g33948, g33949, g33950, g33959, g34201, g34221, g34232, g34233, 
        g34234, g34235, g34236, g34237, g34238, g34239, g34240, g34383, g34425, 
        g34435, g34436, g34437, g34597, g34788, g34839, g34913, g34915, g34917, 
        g34919, g34921, g34923, g34925, g34927, g34956, g34972, test_se, 
        test_si );

    always // clock with period 1000ns
    begin
        clk = 1;
        #500;
        clk = !clk;
        #500;
    end
    


    // Test Patterns
    initial 
    begin

        // Create a file for writing the outputs of the testbench
        file = $fopen("tb_s38584.txt", "w");

        // Flash the reset on the DUT
        rst = 1;
        #1000;
        rst = 0;

        for (i=0; i < 12; i = i+1)
        begin

            // Have the first test be non random.
            if (i < 2)

                // First index, test all ones
                if (i==0)
                begin

                    // assign all 1's to the inputs
                    g35 = 1;
                    g36 = 1;
                    g6744 = 1;
                    g6745 = 1;
                    g6746 = 1;
                    g6747 = 1;
                    g6748 = 1;
                    g6749 = 1;
                    g6750 = 1;
                    g6751 = 1;
                    g6752 = 1;
                    g6753 = 1;
                    test_se = 1;
                    test_si = 1;
                end

                // Second index, test all zeros
                else
                begin

                    // assign all 0's to the inputs
                    g35 = 0;
                    g36 = 0;
                    g6744 = 0;
                    g6745 = 0;
                    g6746 = 0;
                    g6747 = 0;
                    g6748 = 0;
                    g6749 = 0;
                    g6750 = 0;
                    g6751 = 0;
                    g6752 = 0;
                    g6753 = 0;
                    test_se = 0; 
                    test_si = 0;
                end

            else
            begin
                // assign random data
                {g35, g36, g6744, g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6752, g6753, test_se, test_si} = $random;
            end
            
            // write to the file 
            $fwrite(file,"Input Pattern: %b\n", {g35, g36, g6744, g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6752, g6753, test_se, test_si});
            $fwrite(file,"Output Pattern: %b\n", {g7243, g7245, g7257, g7260, g7540, g7916, g7946, g8132, g8178, g8215,
                                                    g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353, g8358, g8398,
                                                    g8403, g8416, g8475, g8719, g8783, g8784, g8785, g8786, g8787, g8788,
                                                    g8789, g8839, g8870, g8915, g8916, g8917, g8918, g8919, g8920, g9019,
                                                    g9048, g9251, g9497, g9553, g9555, g9615, g9617, g9680, g9682, g9741,
                                                    g9743, g9817, g10122, g10306, g10500, g10527, g11349, g11388, g11418,
                                                    g11447, g11678, g11770, g12184, g12238, g12300, g12350, g12368,
                                                    g12422, g12470, g12832, g12919, g12923, g13039, g13049, g13068,
                                                    g13085, g13099, g13259, g13272, g13865, g13881, g13895, g13906,
                                                    g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201,
                                                    g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673,
                                                    g14694, g14705, g14738, g14749, g14779, g14828, g16603, g16624,
                                                    g16627, g16656, g16659, g16686, g16693, g16718, g16722, g16744,
                                                    g16748, g16775, g16874, g16924, g16955, g17291, g17316, g17320,
                                                    g17400, g17404, g17423, g17519, g17577, g17580, g17604, g17607,
                                                    g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711,
                                                    g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787,
                                                    g17813, g17819, g17845, g17871, g18092, g18094, g18095, g18096,
                                                    g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357,
                                                    g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176,
                                                    g21245, g21270, g21292, g21698, g21727, g23002, g23190, g23612,
                                                    g23652, g23683, g23759, g24151, g25114, g25167, g25219, g25259,
                                                    g25582, g25583, g25584, g25585, g25586, g25587, g25588, g25589,
                                                    g25590, g26801, g26875, g26876, g26877, g27831, g28030, g28041,
                                                    g28042, g28753, g29210, g29211, g29212, g29213, g29214, g29215,
                                                    g29216, g29217, g29218, g29219, g29220, g29221, g30327, g30329,
                                                    g30330, g30331, g30332, g31521, g31656, g31665, g31793, g31860,
                                                    g31861, g31862, g31863, g32185, g32429, g32454, g32975, g33079,
                                                    g33435, g33533, g33636, g33659, g33874, g33894, g33935, g33945,
                                                    g33946, g33947, g33948, g33949, g33950, g33959, g34201, g34221,
                                                    g34232, g34233, g34234, g34235, g34236, g34237, g34238, g34239,
                                                    g34240, g34383, g34425, g34435, g34436, g34437, g34597, g34788,
                                                    g34839, g34913, g34915, g34917, g34919, g34921, g34923, g34925,
                                                    g34927, g34956, g34972});

            // wait 5000 ns before the next iteration
            #5000;

        end;

    // Close the file
    $fclose(file);
    $finish;
    end

endmodule