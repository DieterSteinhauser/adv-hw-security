VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS

USEMINSPACING OBS ON ;
USEMINSPACING PIN OFF ;
CLEARANCEMEASURE EUCLIDEAN ;


MANUFACTURINGGRID 0.005 ;

MACRO XOR2X1
  CLASS  CORE ;
  FOREIGN XOR2X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.260 BY 7.920 ;
  SYMMETRY X Y  ;
  SITE CORE ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.090 3.430 4.490 3.880 ;
        RECT 4.090 3.480 5.120 3.880 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 0.980 2.530 1.380 2.930 ;
        RECT 5.620 3.480 6.020 3.880 ;
        RECT 5.620 2.630 5.920 3.880 ;
        RECT 5.460 2.630 5.920 3.120 ;
        RECT 0.980 2.630 5.920 2.930 ;
    END
  END B
  PIN GRND
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 1.280 -0.540 1.680 1.490 ;
        RECT 0.000 -0.540 7.260 0.540 ;
        RECT 6.000 -0.540 6.400 1.490 ;
        RECT 3.460 -0.540 3.860 1.900 ;
        RECT 3.440 -0.540 3.860 0.650 ;
    END
  END GRND
  PIN Y
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 4.240 1.250 4.640 2.090 ;
        RECT 6.320 2.110 7.080 2.510 ;
        RECT 5.020 4.280 6.620 4.580 ;
        RECT 6.320 1.790 6.620 4.580 ;
        RECT 4.240 1.790 6.620 2.090 ;
        RECT 5.020 4.280 5.420 6.280 ;
        RECT 4.440 0.840 4.840 1.490 ;
    END
  END Y
  PIN POWR
    DIRECTION INPUT ;
    PORT
      LAYER Metal1 ;
        RECT 2.060 4.070 2.460 8.460 ;
        RECT 0.000 7.380 7.260 8.460 ;
        RECT 3.460 4.280 3.860 8.460 ;
        RECT 0.840 7.270 2.840 8.460 ;
    END
  END POWR
  OBS 
      LAYER Metal1 ;
        RECT 1.280 4.070 1.680 6.670 ;
        RECT 0.500 0.840 0.900 2.090 ;
        RECT 2.060 0.840 2.460 2.090 ;
        RECT 0.380 1.790 3.060 2.090 ;
        RECT 2.660 1.790 3.060 2.290 ;
        RECT 0.380 1.790 0.680 3.770 ;
        RECT 0.380 3.470 3.790 3.770 ;
        RECT 3.390 3.470 3.790 3.880 ;
        RECT 0.500 3.470 0.900 6.670 ;
        RECT 5.220 0.840 5.620 1.490 ;
        RECT 4.240 4.280 4.640 7.080 ;
        RECT 5.800 5.080 6.200 7.080 ;
        RECT 4.240 6.680 6.200 7.080 ;
  END 
END XOR2X1

END LIBRARY
